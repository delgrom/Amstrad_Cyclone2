-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"d4080b0b",
    10 => x"0bbdd808",
    11 => x"0b0b0bbd",
    12 => x"dc080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bddc0c0b",
    16 => x"0b0bbdd8",
    17 => x"0c0b0b0b",
    18 => x"bdd40c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb284",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bdd47080",
    57 => x"c884278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188e304",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbde40c",
    65 => x"9f0bbde8",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bde808ff",
    69 => x"05bde80c",
    70 => x"bde80880",
    71 => x"25eb38bd",
    72 => x"e408ff05",
    73 => x"bde40cbd",
    74 => x"e4088025",
    75 => x"d738800b",
    76 => x"bde80c80",
    77 => x"0bbde40c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbde408",
    97 => x"258f3882",
    98 => x"bd2dbde4",
    99 => x"08ff05bd",
   100 => x"e40c82ff",
   101 => x"04bde408",
   102 => x"bde80853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bde408a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bde8",
   111 => x"088105bd",
   112 => x"e80cbde8",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbde80c",
   116 => x"bde40881",
   117 => x"05bde40c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bd",
   122 => x"e8088105",
   123 => x"bde80cbd",
   124 => x"e808a02e",
   125 => x"0981068e",
   126 => x"38800bbd",
   127 => x"e80cbde4",
   128 => x"088105bd",
   129 => x"e40c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbdec",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbdec0c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bd",
   169 => x"ec088407",
   170 => x"bdec0c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb8e4",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bdec0852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bdd40c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402d0",
   222 => x"050d7d54",
   223 => x"807453bd",
   224 => x"f0525ba9",
   225 => x"a32dbdd4",
   226 => x"087b2e81",
   227 => x"af38bdf4",
   228 => x"0870f80c",
   229 => x"891580f5",
   230 => x"2d8a1680",
   231 => x"f52d7182",
   232 => x"80290588",
   233 => x"1780f52d",
   234 => x"70848080",
   235 => x"2912f40c",
   236 => x"57555658",
   237 => x"a40bec0c",
   238 => x"7aff1958",
   239 => x"5a767b2e",
   240 => x"8b38811a",
   241 => x"77812a58",
   242 => x"5a76f738",
   243 => x"f71a5a81",
   244 => x"5b807825",
   245 => x"80e63879",
   246 => x"52765184",
   247 => x"8b2dbebc",
   248 => x"52bdf051",
   249 => x"abe22dbd",
   250 => x"d408802e",
   251 => x"b838bebc",
   252 => x"5c83fc59",
   253 => x"7b708405",
   254 => x"5d087081",
   255 => x"ff067188",
   256 => x"2a7081ff",
   257 => x"0673902a",
   258 => x"7081ff06",
   259 => x"75982ae8",
   260 => x"0ce80c58",
   261 => x"e80c57e8",
   262 => x"0cfc1a5a",
   263 => x"53788025",
   264 => x"d33888ac",
   265 => x"04bdd408",
   266 => x"5b848058",
   267 => x"bdf051ab",
   268 => x"b42dfc80",
   269 => x"18811858",
   270 => x"5887d104",
   271 => x"86b72d84",
   272 => x"0bec0c7a",
   273 => x"802e8d38",
   274 => x"b8e85191",
   275 => x"c92d8fcc",
   276 => x"2d88da04",
   277 => x"bba45191",
   278 => x"c92d7abd",
   279 => x"d40c02b0",
   280 => x"050d0402",
   281 => x"d4050d80",
   282 => x"55840bec",
   283 => x"0c8fad2d",
   284 => x"8c972d81",
   285 => x"f82da098",
   286 => x"2dbdd408",
   287 => x"752e8382",
   288 => x"388c0bec",
   289 => x"0cb7a452",
   290 => x"bdf051a9",
   291 => x"a32dbdd4",
   292 => x"08752e81",
   293 => x"8338bdf4",
   294 => x"0875ff12",
   295 => x"595b5876",
   296 => x"752e8b38",
   297 => x"811a7781",
   298 => x"2a585a76",
   299 => x"f738f71a",
   300 => x"5a807825",
   301 => x"80e23879",
   302 => x"52765184",
   303 => x"8b2dbebc",
   304 => x"52bdf051",
   305 => x"abe22dbd",
   306 => x"d408802e",
   307 => x"b838bebc",
   308 => x"5b83fc59",
   309 => x"7a708405",
   310 => x"5c087081",
   311 => x"ff067188",
   312 => x"2a7081ff",
   313 => x"0673902a",
   314 => x"7081ff06",
   315 => x"75982ae8",
   316 => x"0ce80c58",
   317 => x"e80c57e8",
   318 => x"0cfc1a5a",
   319 => x"53788025",
   320 => x"d3388a88",
   321 => x"04848058",
   322 => x"bdf051ab",
   323 => x"b42dfc80",
   324 => x"18811858",
   325 => x"5889b104",
   326 => x"bdf408f8",
   327 => x"0c86b72d",
   328 => x"840bec0c",
   329 => x"86f651b1",
   330 => x"fc2db8e8",
   331 => x"5191c92d",
   332 => x"8fcc2d8c",
   333 => x"a32d91d9",
   334 => x"2db9880b",
   335 => x"80f52d70",
   336 => x"822b9c06",
   337 => x"b8fc0b80",
   338 => x"f52d8306",
   339 => x"7107b994",
   340 => x"0b80f52d",
   341 => x"70852ba0",
   342 => x"06b9a00b",
   343 => x"80f52d70",
   344 => x"862b80c0",
   345 => x"06747307",
   346 => x"07b9ac0b",
   347 => x"80f52d70",
   348 => x"872b8180",
   349 => x"06b9b80b",
   350 => x"80f52d70",
   351 => x"882b8280",
   352 => x"06747307",
   353 => x"07b9c40b",
   354 => x"80f52d70",
   355 => x"892b8480",
   356 => x"06b9d00b",
   357 => x"80f52d70",
   358 => x"8a2b8880",
   359 => x"06747307",
   360 => x"07b9dc0b",
   361 => x"80f52d70",
   362 => x"8b2b9080",
   363 => x"06b9e80b",
   364 => x"80f52d70",
   365 => x"8c2ba080",
   366 => x"06747307",
   367 => x"07b9f40b",
   368 => x"80f52d70",
   369 => x"8d2b81c0",
   370 => x"8006ba80",
   371 => x"0b80f52d",
   372 => x"708f2b82",
   373 => x"80800674",
   374 => x"730707fc",
   375 => x"0c545454",
   376 => x"54545454",
   377 => x"54545454",
   378 => x"54545454",
   379 => x"545b5452",
   380 => x"57545486",
   381 => x"53bdd408",
   382 => x"83388453",
   383 => x"72ec0c8a",
   384 => x"b304800b",
   385 => x"bdd40c02",
   386 => x"ac050d04",
   387 => x"71980c04",
   388 => x"ffb008bd",
   389 => x"d40c0481",
   390 => x"0bffb00c",
   391 => x"04800bff",
   392 => x"b00c0402",
   393 => x"f4050d8d",
   394 => x"a504bdd4",
   395 => x"0881f02e",
   396 => x"09810689",
   397 => x"38810bbc",
   398 => x"880c8da5",
   399 => x"04bdd408",
   400 => x"81e02e09",
   401 => x"81068938",
   402 => x"810bbc8c",
   403 => x"0c8da504",
   404 => x"bdd40852",
   405 => x"bc8c0880",
   406 => x"2e8838bd",
   407 => x"d4088180",
   408 => x"05527184",
   409 => x"2c728f06",
   410 => x"5353bc88",
   411 => x"08802e99",
   412 => x"38728429",
   413 => x"bbc80572",
   414 => x"1381712b",
   415 => x"70097308",
   416 => x"06730c51",
   417 => x"53538d9b",
   418 => x"04728429",
   419 => x"bbc80572",
   420 => x"1383712b",
   421 => x"72080772",
   422 => x"0c535380",
   423 => x"0bbc8c0c",
   424 => x"800bbc88",
   425 => x"0cbdfc51",
   426 => x"8ea62dbd",
   427 => x"d408ff24",
   428 => x"fef83880",
   429 => x"0bbdd40c",
   430 => x"028c050d",
   431 => x"0402f805",
   432 => x"0dbbc852",
   433 => x"8f518072",
   434 => x"70840554",
   435 => x"0cff1151",
   436 => x"708025f2",
   437 => x"38028805",
   438 => x"0d0402f0",
   439 => x"050d7551",
   440 => x"8c9d2d70",
   441 => x"822cfc06",
   442 => x"bbc81172",
   443 => x"109e0671",
   444 => x"0870722a",
   445 => x"70830682",
   446 => x"742b7009",
   447 => x"7406760c",
   448 => x"54515657",
   449 => x"5351538c",
   450 => x"972d71bd",
   451 => x"d40c0290",
   452 => x"050d0402",
   453 => x"fc050d72",
   454 => x"5180710c",
   455 => x"800b8412",
   456 => x"0c028405",
   457 => x"0d0402f0",
   458 => x"050d7570",
   459 => x"08841208",
   460 => x"535353ff",
   461 => x"5471712e",
   462 => x"a8388c9d",
   463 => x"2d841308",
   464 => x"70842914",
   465 => x"88117008",
   466 => x"7081ff06",
   467 => x"84180881",
   468 => x"11870684",
   469 => x"1a0c5351",
   470 => x"55515151",
   471 => x"8c972d71",
   472 => x"5473bdd4",
   473 => x"0c029005",
   474 => x"0d0402f8",
   475 => x"050d8c9d",
   476 => x"2de00870",
   477 => x"8b2a7081",
   478 => x"06515252",
   479 => x"70802e9d",
   480 => x"38bdfc08",
   481 => x"708429be",
   482 => x"84057381",
   483 => x"ff06710c",
   484 => x"5151bdfc",
   485 => x"08811187",
   486 => x"06bdfc0c",
   487 => x"51800bbe",
   488 => x"a40c8c90",
   489 => x"2d8c972d",
   490 => x"0288050d",
   491 => x"0402fc05",
   492 => x"0dbdfc51",
   493 => x"8e932d8d",
   494 => x"bd2d8eea",
   495 => x"518c8c2d",
   496 => x"0284050d",
   497 => x"04bea808",
   498 => x"bdd40c04",
   499 => x"02fc050d",
   500 => x"8fd6048c",
   501 => x"a32d80f6",
   502 => x"518dda2d",
   503 => x"bdd408f3",
   504 => x"3880da51",
   505 => x"8dda2dbd",
   506 => x"d408e838",
   507 => x"bdd408bc",
   508 => x"940cbdd4",
   509 => x"085184f0",
   510 => x"2d028405",
   511 => x"0d0402ec",
   512 => x"050d7654",
   513 => x"8052870b",
   514 => x"881580f5",
   515 => x"2d565374",
   516 => x"72248338",
   517 => x"a0537251",
   518 => x"82f92d81",
   519 => x"128b1580",
   520 => x"f52d5452",
   521 => x"727225de",
   522 => x"38029405",
   523 => x"0d0402f0",
   524 => x"050dbea8",
   525 => x"085481f8",
   526 => x"2d800bbe",
   527 => x"ac0c7308",
   528 => x"802e8180",
   529 => x"38820bbd",
   530 => x"e80cbeac",
   531 => x"088f06bd",
   532 => x"e40c7308",
   533 => x"5271832e",
   534 => x"96387183",
   535 => x"26893871",
   536 => x"812eaf38",
   537 => x"91af0471",
   538 => x"852e9f38",
   539 => x"91af0488",
   540 => x"1480f52d",
   541 => x"841508b7",
   542 => x"b0535452",
   543 => x"85fe2d71",
   544 => x"84291370",
   545 => x"08525291",
   546 => x"b3047351",
   547 => x"8ffe2d91",
   548 => x"af04bc90",
   549 => x"08881508",
   550 => x"2c708106",
   551 => x"51527180",
   552 => x"2e8738b7",
   553 => x"b45191ac",
   554 => x"04b7b851",
   555 => x"85fe2d84",
   556 => x"14085185",
   557 => x"fe2dbeac",
   558 => x"088105be",
   559 => x"ac0c8c14",
   560 => x"5490be04",
   561 => x"0290050d",
   562 => x"0471bea8",
   563 => x"0c90ae2d",
   564 => x"beac08ff",
   565 => x"05beb00c",
   566 => x"0402e805",
   567 => x"0dbea808",
   568 => x"beb40857",
   569 => x"5587518d",
   570 => x"da2dbdd4",
   571 => x"08812a70",
   572 => x"81065152",
   573 => x"71802ea0",
   574 => x"3891ff04",
   575 => x"8ca32d87",
   576 => x"518dda2d",
   577 => x"bdd408f4",
   578 => x"38bc9408",
   579 => x"813270bc",
   580 => x"940c7052",
   581 => x"5284f02d",
   582 => x"80fe518d",
   583 => x"da2dbdd4",
   584 => x"08802ea6",
   585 => x"38bc9408",
   586 => x"802e9138",
   587 => x"800bbc94",
   588 => x"0c805184",
   589 => x"f02d92bc",
   590 => x"048ca32d",
   591 => x"80fe518d",
   592 => x"da2dbdd4",
   593 => x"08f33886",
   594 => x"e22dbc94",
   595 => x"08903881",
   596 => x"fd518dda",
   597 => x"2d81fa51",
   598 => x"8dda2d98",
   599 => x"8f0481f5",
   600 => x"518dda2d",
   601 => x"bdd40881",
   602 => x"2a708106",
   603 => x"51527180",
   604 => x"2eaf38be",
   605 => x"b0085271",
   606 => x"802e8938",
   607 => x"ff12beb0",
   608 => x"0c93a104",
   609 => x"beac0810",
   610 => x"beac0805",
   611 => x"70842916",
   612 => x"51528812",
   613 => x"08802e89",
   614 => x"38ff5188",
   615 => x"12085271",
   616 => x"2d81f251",
   617 => x"8dda2dbd",
   618 => x"d408812a",
   619 => x"70810651",
   620 => x"5271802e",
   621 => x"b138beac",
   622 => x"08ff11be",
   623 => x"b0085653",
   624 => x"53737225",
   625 => x"89388114",
   626 => x"beb00c93",
   627 => x"e6047210",
   628 => x"13708429",
   629 => x"16515288",
   630 => x"1208802e",
   631 => x"8938fe51",
   632 => x"88120852",
   633 => x"712d81fd",
   634 => x"518dda2d",
   635 => x"bdd40881",
   636 => x"2a708106",
   637 => x"51527180",
   638 => x"2ead38be",
   639 => x"b008802e",
   640 => x"8938800b",
   641 => x"beb00c94",
   642 => x"a704beac",
   643 => x"0810beac",
   644 => x"08057084",
   645 => x"29165152",
   646 => x"88120880",
   647 => x"2e8938fd",
   648 => x"51881208",
   649 => x"52712d81",
   650 => x"fa518dda",
   651 => x"2dbdd408",
   652 => x"812a7081",
   653 => x"06515271",
   654 => x"802eae38",
   655 => x"beac08ff",
   656 => x"115452be",
   657 => x"b0087325",
   658 => x"883872be",
   659 => x"b00c94e9",
   660 => x"04711012",
   661 => x"70842916",
   662 => x"51528812",
   663 => x"08802e89",
   664 => x"38fc5188",
   665 => x"12085271",
   666 => x"2dbeb008",
   667 => x"70535473",
   668 => x"802e8a38",
   669 => x"8c15ff15",
   670 => x"555594ef",
   671 => x"04820bbd",
   672 => x"e80c718f",
   673 => x"06bde40c",
   674 => x"81eb518d",
   675 => x"da2dbdd4",
   676 => x"08812a70",
   677 => x"81065152",
   678 => x"71802ead",
   679 => x"38740885",
   680 => x"2e098106",
   681 => x"a4388815",
   682 => x"80f52dff",
   683 => x"05527188",
   684 => x"1681b72d",
   685 => x"71982b52",
   686 => x"71802588",
   687 => x"38800b88",
   688 => x"1681b72d",
   689 => x"74518ffe",
   690 => x"2d81f451",
   691 => x"8dda2dbd",
   692 => x"d408812a",
   693 => x"70810651",
   694 => x"5271802e",
   695 => x"b3387408",
   696 => x"852e0981",
   697 => x"06aa3888",
   698 => x"1580f52d",
   699 => x"81055271",
   700 => x"881681b7",
   701 => x"2d7181ff",
   702 => x"068b1680",
   703 => x"f52d5452",
   704 => x"72722787",
   705 => x"38728816",
   706 => x"81b72d74",
   707 => x"518ffe2d",
   708 => x"80da518d",
   709 => x"da2dbdd4",
   710 => x"08812a70",
   711 => x"81065152",
   712 => x"71802e81",
   713 => x"a638bea8",
   714 => x"08beb008",
   715 => x"55537380",
   716 => x"2e8a388c",
   717 => x"13ff1555",
   718 => x"5396ae04",
   719 => x"72085271",
   720 => x"822ea638",
   721 => x"71822689",
   722 => x"3871812e",
   723 => x"a93897cb",
   724 => x"0471832e",
   725 => x"b1387184",
   726 => x"2e098106",
   727 => x"80ed3888",
   728 => x"13085191",
   729 => x"c92d97cb",
   730 => x"04beb008",
   731 => x"51881308",
   732 => x"52712d97",
   733 => x"cb04810b",
   734 => x"8814082b",
   735 => x"bc900832",
   736 => x"bc900c97",
   737 => x"a1048813",
   738 => x"80f52d81",
   739 => x"058b1480",
   740 => x"f52d5354",
   741 => x"71742483",
   742 => x"38805473",
   743 => x"881481b7",
   744 => x"2d90ae2d",
   745 => x"97cb0475",
   746 => x"08802ea2",
   747 => x"38750851",
   748 => x"8dda2dbd",
   749 => x"d4088106",
   750 => x"5271802e",
   751 => x"8b38beb0",
   752 => x"08518416",
   753 => x"0852712d",
   754 => x"88165675",
   755 => x"da388054",
   756 => x"800bbde8",
   757 => x"0c738f06",
   758 => x"bde40ca0",
   759 => x"5273beb0",
   760 => x"082e0981",
   761 => x"069838be",
   762 => x"ac08ff05",
   763 => x"74327009",
   764 => x"81057072",
   765 => x"079f2a91",
   766 => x"71315151",
   767 => x"53537151",
   768 => x"82f92d81",
   769 => x"14548e74",
   770 => x"25c638bc",
   771 => x"94085271",
   772 => x"bdd40c02",
   773 => x"98050d04",
   774 => x"02f4050d",
   775 => x"d45281ff",
   776 => x"720c7108",
   777 => x"5381ff72",
   778 => x"0c72882b",
   779 => x"83fe8006",
   780 => x"72087081",
   781 => x"ff065152",
   782 => x"5381ff72",
   783 => x"0c727107",
   784 => x"882b7208",
   785 => x"7081ff06",
   786 => x"51525381",
   787 => x"ff720c72",
   788 => x"7107882b",
   789 => x"72087081",
   790 => x"ff067207",
   791 => x"bdd40c52",
   792 => x"53028c05",
   793 => x"0d0402f4",
   794 => x"050d7476",
   795 => x"7181ff06",
   796 => x"d40c5353",
   797 => x"beb80885",
   798 => x"3871892b",
   799 => x"5271982a",
   800 => x"d40c7190",
   801 => x"2a7081ff",
   802 => x"06d40c51",
   803 => x"71882a70",
   804 => x"81ff06d4",
   805 => x"0c517181",
   806 => x"ff06d40c",
   807 => x"72902a70",
   808 => x"81ff06d4",
   809 => x"0c51d408",
   810 => x"7081ff06",
   811 => x"515182b8",
   812 => x"bf527081",
   813 => x"ff2e0981",
   814 => x"06943881",
   815 => x"ff0bd40c",
   816 => x"d4087081",
   817 => x"ff06ff14",
   818 => x"54515171",
   819 => x"e53870bd",
   820 => x"d40c028c",
   821 => x"050d0402",
   822 => x"fc050d81",
   823 => x"c75181ff",
   824 => x"0bd40cff",
   825 => x"11517080",
   826 => x"25f43802",
   827 => x"84050d04",
   828 => x"02f4050d",
   829 => x"81ff0bd4",
   830 => x"0c935380",
   831 => x"5287fc80",
   832 => x"c15198e6",
   833 => x"2dbdd408",
   834 => x"8b3881ff",
   835 => x"0bd40c81",
   836 => x"539a9d04",
   837 => x"99d72dff",
   838 => x"135372df",
   839 => x"3872bdd4",
   840 => x"0c028c05",
   841 => x"0d0402ec",
   842 => x"050d810b",
   843 => x"beb80c84",
   844 => x"54d00870",
   845 => x"8f2a7081",
   846 => x"06515153",
   847 => x"72f33872",
   848 => x"d00c99d7",
   849 => x"2db7bc51",
   850 => x"85fe2dd0",
   851 => x"08708f2a",
   852 => x"70810651",
   853 => x"515372f3",
   854 => x"38810bd0",
   855 => x"0cb15380",
   856 => x"5284d480",
   857 => x"c05198e6",
   858 => x"2dbdd408",
   859 => x"812e9338",
   860 => x"72822ebd",
   861 => x"38ff1353",
   862 => x"72e538ff",
   863 => x"145473ff",
   864 => x"b03899d7",
   865 => x"2d83aa52",
   866 => x"849c80c8",
   867 => x"5198e62d",
   868 => x"bdd40881",
   869 => x"2e098106",
   870 => x"92389898",
   871 => x"2dbdd408",
   872 => x"83ffff06",
   873 => x"537283aa",
   874 => x"2e9d3899",
   875 => x"f02d9bc2",
   876 => x"04b7c851",
   877 => x"85fe2d80",
   878 => x"539d9004",
   879 => x"b7e05185",
   880 => x"fe2d8054",
   881 => x"9ce20481",
   882 => x"ff0bd40c",
   883 => x"b15499d7",
   884 => x"2d8fcf53",
   885 => x"805287fc",
   886 => x"80f75198",
   887 => x"e62dbdd4",
   888 => x"0855bdd4",
   889 => x"08812e09",
   890 => x"81069b38",
   891 => x"81ff0bd4",
   892 => x"0c820a52",
   893 => x"849c80e9",
   894 => x"5198e62d",
   895 => x"bdd40880",
   896 => x"2e8d3899",
   897 => x"d72dff13",
   898 => x"5372c938",
   899 => x"9cd50481",
   900 => x"ff0bd40c",
   901 => x"bdd40852",
   902 => x"87fc80fa",
   903 => x"5198e62d",
   904 => x"bdd408b1",
   905 => x"3881ff0b",
   906 => x"d40cd408",
   907 => x"5381ff0b",
   908 => x"d40c81ff",
   909 => x"0bd40c81",
   910 => x"ff0bd40c",
   911 => x"81ff0bd4",
   912 => x"0c72862a",
   913 => x"70810676",
   914 => x"56515372",
   915 => x"9538bdd4",
   916 => x"08549ce2",
   917 => x"0473822e",
   918 => x"fee238ff",
   919 => x"145473fe",
   920 => x"ed3873be",
   921 => x"b80c738b",
   922 => x"38815287",
   923 => x"fc80d051",
   924 => x"98e62d81",
   925 => x"ff0bd40c",
   926 => x"d008708f",
   927 => x"2a708106",
   928 => x"51515372",
   929 => x"f33872d0",
   930 => x"0c81ff0b",
   931 => x"d40c8153",
   932 => x"72bdd40c",
   933 => x"0294050d",
   934 => x"0402e805",
   935 => x"0d785580",
   936 => x"5681ff0b",
   937 => x"d40cd008",
   938 => x"708f2a70",
   939 => x"81065151",
   940 => x"5372f338",
   941 => x"82810bd0",
   942 => x"0c81ff0b",
   943 => x"d40c7752",
   944 => x"87fc80d1",
   945 => x"5198e62d",
   946 => x"80dbc6df",
   947 => x"54bdd408",
   948 => x"802e8a38",
   949 => x"b8805185",
   950 => x"fe2d9eb0",
   951 => x"0481ff0b",
   952 => x"d40cd408",
   953 => x"7081ff06",
   954 => x"51537281",
   955 => x"fe2e0981",
   956 => x"069d3880",
   957 => x"ff539898",
   958 => x"2dbdd408",
   959 => x"75708405",
   960 => x"570cff13",
   961 => x"53728025",
   962 => x"ed388156",
   963 => x"9e9504ff",
   964 => x"145473c9",
   965 => x"3881ff0b",
   966 => x"d40c81ff",
   967 => x"0bd40cd0",
   968 => x"08708f2a",
   969 => x"70810651",
   970 => x"515372f3",
   971 => x"3872d00c",
   972 => x"75bdd40c",
   973 => x"0298050d",
   974 => x"0402e805",
   975 => x"0d77797b",
   976 => x"58555580",
   977 => x"53727625",
   978 => x"a3387470",
   979 => x"81055680",
   980 => x"f52d7470",
   981 => x"81055680",
   982 => x"f52d5252",
   983 => x"71712e86",
   984 => x"3881519e",
   985 => x"ee048113",
   986 => x"539ec504",
   987 => x"805170bd",
   988 => x"d40c0298",
   989 => x"050d0402",
   990 => x"ec050d76",
   991 => x"5574802e",
   992 => x"be389a15",
   993 => x"80e02d51",
   994 => x"acbb2dbd",
   995 => x"d408bdd4",
   996 => x"0880c4ec",
   997 => x"0cbdd408",
   998 => x"545480c4",
   999 => x"c808802e",
  1000 => x"99389415",
  1001 => x"80e02d51",
  1002 => x"acbb2dbd",
  1003 => x"d408902b",
  1004 => x"83fff00a",
  1005 => x"06707507",
  1006 => x"51537280",
  1007 => x"c4ec0c80",
  1008 => x"c4ec0853",
  1009 => x"72802e9d",
  1010 => x"3880c4c0",
  1011 => x"08fe1471",
  1012 => x"2980c4d4",
  1013 => x"080580c4",
  1014 => x"f00c7084",
  1015 => x"2b80c4cc",
  1016 => x"0c54a093",
  1017 => x"0480c4d8",
  1018 => x"0880c4ec",
  1019 => x"0c80c4dc",
  1020 => x"0880c4f0",
  1021 => x"0c80c4c8",
  1022 => x"08802e8b",
  1023 => x"3880c4c0",
  1024 => x"08842b53",
  1025 => x"a08e0480",
  1026 => x"c4e00884",
  1027 => x"2b537280",
  1028 => x"c4cc0c02",
  1029 => x"94050d04",
  1030 => x"02d8050d",
  1031 => x"800b80c4",
  1032 => x"c80c8454",
  1033 => x"9aa62dbd",
  1034 => x"d408802e",
  1035 => x"9538bebc",
  1036 => x"5280519d",
  1037 => x"992dbdd4",
  1038 => x"08802e86",
  1039 => x"38fe54a0",
  1040 => x"ca04ff14",
  1041 => x"54738024",
  1042 => x"db38738c",
  1043 => x"38b89051",
  1044 => x"85fe2d73",
  1045 => x"55a5f404",
  1046 => x"8056810b",
  1047 => x"80c4f40c",
  1048 => x"8853b8a4",
  1049 => x"52bef251",
  1050 => x"9eb92dbd",
  1051 => x"d408762e",
  1052 => x"09810688",
  1053 => x"38bdd408",
  1054 => x"80c4f40c",
  1055 => x"8853b8b0",
  1056 => x"52bf8e51",
  1057 => x"9eb92dbd",
  1058 => x"d4088838",
  1059 => x"bdd40880",
  1060 => x"c4f40c80",
  1061 => x"c4f40880",
  1062 => x"2e80fc38",
  1063 => x"80c2820b",
  1064 => x"80f52d80",
  1065 => x"c2830b80",
  1066 => x"f52d7198",
  1067 => x"2b71902b",
  1068 => x"0780c284",
  1069 => x"0b80f52d",
  1070 => x"70882b72",
  1071 => x"0780c285",
  1072 => x"0b80f52d",
  1073 => x"710780c2",
  1074 => x"ba0b80f5",
  1075 => x"2d80c2bb",
  1076 => x"0b80f52d",
  1077 => x"71882b07",
  1078 => x"535f5452",
  1079 => x"5a565755",
  1080 => x"7381abaa",
  1081 => x"2e098106",
  1082 => x"8d387551",
  1083 => x"ac8b2dbd",
  1084 => x"d40856a2",
  1085 => x"83047382",
  1086 => x"d4d52e87",
  1087 => x"38b8bc51",
  1088 => x"a2c504be",
  1089 => x"bc527551",
  1090 => x"9d992dbd",
  1091 => x"d40855bd",
  1092 => x"d408802e",
  1093 => x"83de3888",
  1094 => x"53b8b052",
  1095 => x"bf8e519e",
  1096 => x"b92dbdd4",
  1097 => x"088a3881",
  1098 => x"0b80c4c8",
  1099 => x"0ca2cb04",
  1100 => x"8853b8a4",
  1101 => x"52bef251",
  1102 => x"9eb92dbd",
  1103 => x"d408802e",
  1104 => x"8a38b8d0",
  1105 => x"5185fe2d",
  1106 => x"a3a70480",
  1107 => x"c2ba0b80",
  1108 => x"f52d5473",
  1109 => x"80d52e09",
  1110 => x"810680cb",
  1111 => x"3880c2bb",
  1112 => x"0b80f52d",
  1113 => x"547381aa",
  1114 => x"2e098106",
  1115 => x"ba38800b",
  1116 => x"bebc0b80",
  1117 => x"f52d5654",
  1118 => x"7481e92e",
  1119 => x"83388154",
  1120 => x"7481eb2e",
  1121 => x"8c388055",
  1122 => x"73752e09",
  1123 => x"810682e4",
  1124 => x"38bec70b",
  1125 => x"80f52d55",
  1126 => x"748d38be",
  1127 => x"c80b80f5",
  1128 => x"2d547382",
  1129 => x"2e863880",
  1130 => x"55a5f404",
  1131 => x"bec90b80",
  1132 => x"f52d7080",
  1133 => x"c4c00cff",
  1134 => x"0580c4c4",
  1135 => x"0cbeca0b",
  1136 => x"80f52dbe",
  1137 => x"cb0b80f5",
  1138 => x"2d587605",
  1139 => x"77828029",
  1140 => x"057080c4",
  1141 => x"d00cbecc",
  1142 => x"0b80f52d",
  1143 => x"7080c4e4",
  1144 => x"0c80c4c8",
  1145 => x"08595758",
  1146 => x"76802e81",
  1147 => x"ac388853",
  1148 => x"b8b052bf",
  1149 => x"8e519eb9",
  1150 => x"2dbdd408",
  1151 => x"81f63880",
  1152 => x"c4c00870",
  1153 => x"842b80c4",
  1154 => x"cc0c7080",
  1155 => x"c4e00cbe",
  1156 => x"e10b80f5",
  1157 => x"2dbee00b",
  1158 => x"80f52d71",
  1159 => x"82802905",
  1160 => x"bee20b80",
  1161 => x"f52d7084",
  1162 => x"80802912",
  1163 => x"bee30b80",
  1164 => x"f52d7081",
  1165 => x"800a2912",
  1166 => x"7080c4e8",
  1167 => x"0c80c4e4",
  1168 => x"08712980",
  1169 => x"c4d00805",
  1170 => x"7080c4d4",
  1171 => x"0cbee90b",
  1172 => x"80f52dbe",
  1173 => x"e80b80f5",
  1174 => x"2d718280",
  1175 => x"2905beea",
  1176 => x"0b80f52d",
  1177 => x"70848080",
  1178 => x"2912beeb",
  1179 => x"0b80f52d",
  1180 => x"70982b81",
  1181 => x"f00a0672",
  1182 => x"057080c4",
  1183 => x"d80cfe11",
  1184 => x"7e297705",
  1185 => x"80c4dc0c",
  1186 => x"52595243",
  1187 => x"545e5152",
  1188 => x"59525d57",
  1189 => x"5957a5ed",
  1190 => x"04bece0b",
  1191 => x"80f52dbe",
  1192 => x"cd0b80f5",
  1193 => x"2d718280",
  1194 => x"29057080",
  1195 => x"c4cc0c70",
  1196 => x"a02983ff",
  1197 => x"0570892a",
  1198 => x"7080c4e0",
  1199 => x"0cbed30b",
  1200 => x"80f52dbe",
  1201 => x"d20b80f5",
  1202 => x"2d718280",
  1203 => x"29057080",
  1204 => x"c4e80c7b",
  1205 => x"71291e70",
  1206 => x"80c4dc0c",
  1207 => x"7d80c4d8",
  1208 => x"0c730580",
  1209 => x"c4d40c55",
  1210 => x"5e515155",
  1211 => x"5580519e",
  1212 => x"f72d8155",
  1213 => x"74bdd40c",
  1214 => x"02a8050d",
  1215 => x"0402ec05",
  1216 => x"0d767087",
  1217 => x"2c7180ff",
  1218 => x"06555654",
  1219 => x"80c4c808",
  1220 => x"8a387388",
  1221 => x"2c7481ff",
  1222 => x"065455be",
  1223 => x"bc5280c4",
  1224 => x"d0081551",
  1225 => x"9d992dbd",
  1226 => x"d40854bd",
  1227 => x"d408802e",
  1228 => x"b43880c4",
  1229 => x"c808802e",
  1230 => x"98387284",
  1231 => x"29bebc05",
  1232 => x"70085253",
  1233 => x"ac8b2dbd",
  1234 => x"d408f00a",
  1235 => x"0653a6e3",
  1236 => x"047210be",
  1237 => x"bc057080",
  1238 => x"e02d5253",
  1239 => x"acbb2dbd",
  1240 => x"d4085372",
  1241 => x"5473bdd4",
  1242 => x"0c029405",
  1243 => x"0d0402e0",
  1244 => x"050d7970",
  1245 => x"842c80c4",
  1246 => x"f0080571",
  1247 => x"8f065255",
  1248 => x"53728938",
  1249 => x"bebc5273",
  1250 => x"519d992d",
  1251 => x"72a029be",
  1252 => x"bc055480",
  1253 => x"7480f52d",
  1254 => x"56537473",
  1255 => x"2e833881",
  1256 => x"537481e5",
  1257 => x"2e81f138",
  1258 => x"81707406",
  1259 => x"54587280",
  1260 => x"2e81e538",
  1261 => x"8b1480f5",
  1262 => x"2d70832a",
  1263 => x"79065856",
  1264 => x"769938bc",
  1265 => x"98085372",
  1266 => x"89387280",
  1267 => x"c2bc0b81",
  1268 => x"b72d76bc",
  1269 => x"980c7353",
  1270 => x"a99a0475",
  1271 => x"8f2e0981",
  1272 => x"0681b538",
  1273 => x"749f068d",
  1274 => x"2980c2af",
  1275 => x"11515381",
  1276 => x"1480f52d",
  1277 => x"73708105",
  1278 => x"5581b72d",
  1279 => x"831480f5",
  1280 => x"2d737081",
  1281 => x"055581b7",
  1282 => x"2d851480",
  1283 => x"f52d7370",
  1284 => x"81055581",
  1285 => x"b72d8714",
  1286 => x"80f52d73",
  1287 => x"70810555",
  1288 => x"81b72d89",
  1289 => x"1480f52d",
  1290 => x"73708105",
  1291 => x"5581b72d",
  1292 => x"8e1480f5",
  1293 => x"2d737081",
  1294 => x"055581b7",
  1295 => x"2d901480",
  1296 => x"f52d7370",
  1297 => x"81055581",
  1298 => x"b72d9214",
  1299 => x"80f52d73",
  1300 => x"70810555",
  1301 => x"81b72d94",
  1302 => x"1480f52d",
  1303 => x"73708105",
  1304 => x"5581b72d",
  1305 => x"961480f5",
  1306 => x"2d737081",
  1307 => x"055581b7",
  1308 => x"2d981480",
  1309 => x"f52d7370",
  1310 => x"81055581",
  1311 => x"b72d9c14",
  1312 => x"80f52d73",
  1313 => x"70810555",
  1314 => x"81b72d9e",
  1315 => x"1480f52d",
  1316 => x"7381b72d",
  1317 => x"77bc980c",
  1318 => x"805372bd",
  1319 => x"d40c02a0",
  1320 => x"050d0402",
  1321 => x"cc050d7e",
  1322 => x"605e5a80",
  1323 => x"0b80c4ec",
  1324 => x"0880c4f0",
  1325 => x"08595c56",
  1326 => x"805880c4",
  1327 => x"cc08782e",
  1328 => x"81b03877",
  1329 => x"8f06a017",
  1330 => x"5754738f",
  1331 => x"38bebc52",
  1332 => x"76518117",
  1333 => x"579d992d",
  1334 => x"bebc5680",
  1335 => x"7680f52d",
  1336 => x"56547474",
  1337 => x"2e833881",
  1338 => x"547481e5",
  1339 => x"2e80f738",
  1340 => x"81707506",
  1341 => x"555c7380",
  1342 => x"2e80eb38",
  1343 => x"8b1680f5",
  1344 => x"2d980659",
  1345 => x"7880df38",
  1346 => x"8b537c52",
  1347 => x"75519eb9",
  1348 => x"2dbdd408",
  1349 => x"80d0389c",
  1350 => x"160851ac",
  1351 => x"8b2dbdd4",
  1352 => x"08841b0c",
  1353 => x"9a1680e0",
  1354 => x"2d51acbb",
  1355 => x"2dbdd408",
  1356 => x"bdd40888",
  1357 => x"1c0cbdd4",
  1358 => x"08555580",
  1359 => x"c4c80880",
  1360 => x"2e983894",
  1361 => x"1680e02d",
  1362 => x"51acbb2d",
  1363 => x"bdd40890",
  1364 => x"2b83fff0",
  1365 => x"0a067016",
  1366 => x"51547388",
  1367 => x"1b0c787a",
  1368 => x"0c7b54ab",
  1369 => x"ab048118",
  1370 => x"5880c4cc",
  1371 => x"087826fe",
  1372 => x"d23880c4",
  1373 => x"c808802e",
  1374 => x"b0387a51",
  1375 => x"a5fd2dbd",
  1376 => x"d408bdd4",
  1377 => x"0880ffff",
  1378 => x"fff80655",
  1379 => x"5b7380ff",
  1380 => x"fffff82e",
  1381 => x"9438bdd4",
  1382 => x"08fe0580",
  1383 => x"c4c00829",
  1384 => x"80c4d408",
  1385 => x"0557a9b8",
  1386 => x"04805473",
  1387 => x"bdd40c02",
  1388 => x"b4050d04",
  1389 => x"02f4050d",
  1390 => x"74700881",
  1391 => x"05710c70",
  1392 => x"0880c4c4",
  1393 => x"08065353",
  1394 => x"718e3888",
  1395 => x"130851a5",
  1396 => x"fd2dbdd4",
  1397 => x"0888140c",
  1398 => x"810bbdd4",
  1399 => x"0c028c05",
  1400 => x"0d0402f0",
  1401 => x"050d7588",
  1402 => x"1108fe05",
  1403 => x"80c4c008",
  1404 => x"2980c4d4",
  1405 => x"08117208",
  1406 => x"80c4c408",
  1407 => x"06057955",
  1408 => x"5354549d",
  1409 => x"992d0290",
  1410 => x"050d0402",
  1411 => x"f4050d74",
  1412 => x"70882a83",
  1413 => x"fe800670",
  1414 => x"72982a07",
  1415 => x"72882b87",
  1416 => x"fc808006",
  1417 => x"73982b81",
  1418 => x"f00a0671",
  1419 => x"730707bd",
  1420 => x"d40c5651",
  1421 => x"5351028c",
  1422 => x"050d0402",
  1423 => x"f8050d02",
  1424 => x"8e0580f5",
  1425 => x"2d74882b",
  1426 => x"077083ff",
  1427 => x"ff06bdd4",
  1428 => x"0c510288",
  1429 => x"050d0402",
  1430 => x"f4050d74",
  1431 => x"76785354",
  1432 => x"52807125",
  1433 => x"97387270",
  1434 => x"81055480",
  1435 => x"f52d7270",
  1436 => x"81055481",
  1437 => x"b72dff11",
  1438 => x"5170eb38",
  1439 => x"807281b7",
  1440 => x"2d028c05",
  1441 => x"0d0402e8",
  1442 => x"050d7756",
  1443 => x"80705654",
  1444 => x"737624b3",
  1445 => x"3880c4cc",
  1446 => x"08742eab",
  1447 => x"387351a6",
  1448 => x"ee2dbdd4",
  1449 => x"08bdd408",
  1450 => x"09810570",
  1451 => x"bdd40807",
  1452 => x"9f2a7705",
  1453 => x"81175757",
  1454 => x"53537476",
  1455 => x"24893880",
  1456 => x"c4cc0874",
  1457 => x"26d73872",
  1458 => x"bdd40c02",
  1459 => x"98050d04",
  1460 => x"02f0050d",
  1461 => x"bdd00816",
  1462 => x"51ad862d",
  1463 => x"bdd40880",
  1464 => x"2e9e388b",
  1465 => x"53bdd408",
  1466 => x"5280c2bc",
  1467 => x"51acd72d",
  1468 => x"80c4f808",
  1469 => x"5473802e",
  1470 => x"873880c2",
  1471 => x"bc51732d",
  1472 => x"0290050d",
  1473 => x"0402dc05",
  1474 => x"0d80705a",
  1475 => x"5574bdd0",
  1476 => x"0825b138",
  1477 => x"80c4cc08",
  1478 => x"752ea938",
  1479 => x"7851a6ee",
  1480 => x"2dbdd408",
  1481 => x"09810570",
  1482 => x"bdd40807",
  1483 => x"9f2a7605",
  1484 => x"811b5b56",
  1485 => x"5474bdd0",
  1486 => x"08258938",
  1487 => x"80c4cc08",
  1488 => x"7926d938",
  1489 => x"80557880",
  1490 => x"c4cc0827",
  1491 => x"81d43878",
  1492 => x"51a6ee2d",
  1493 => x"bdd40880",
  1494 => x"2e81a838",
  1495 => x"bdd4088b",
  1496 => x"0580f52d",
  1497 => x"70842a70",
  1498 => x"81067710",
  1499 => x"78842b80",
  1500 => x"c2bc0b80",
  1501 => x"f52d5c5c",
  1502 => x"53515556",
  1503 => x"73802e80",
  1504 => x"c9387416",
  1505 => x"822bb0c6",
  1506 => x"0bbca412",
  1507 => x"0c547775",
  1508 => x"311080c4",
  1509 => x"fc115556",
  1510 => x"90747081",
  1511 => x"055681b7",
  1512 => x"2da07481",
  1513 => x"b72d7681",
  1514 => x"ff068116",
  1515 => x"58547380",
  1516 => x"2e8a389c",
  1517 => x"5380c2bc",
  1518 => x"52afc204",
  1519 => x"8b53bdd4",
  1520 => x"085280c4",
  1521 => x"fe1651af",
  1522 => x"fb047416",
  1523 => x"822badd0",
  1524 => x"0bbca412",
  1525 => x"0c547681",
  1526 => x"ff068116",
  1527 => x"58547380",
  1528 => x"2e8a389c",
  1529 => x"5380c2bc",
  1530 => x"52aff204",
  1531 => x"8b53bdd4",
  1532 => x"08527775",
  1533 => x"311080c4",
  1534 => x"fc055176",
  1535 => x"55acd72d",
  1536 => x"b0970474",
  1537 => x"90297531",
  1538 => x"701080c4",
  1539 => x"fc055154",
  1540 => x"bdd40874",
  1541 => x"81b72d81",
  1542 => x"1959748b",
  1543 => x"24a338ae",
  1544 => x"c6047490",
  1545 => x"29753170",
  1546 => x"1080c4fc",
  1547 => x"058c7731",
  1548 => x"57515480",
  1549 => x"7481b72d",
  1550 => x"9e14ff16",
  1551 => x"565474f3",
  1552 => x"3802a405",
  1553 => x"0d0402fc",
  1554 => x"050dbdd0",
  1555 => x"081351ad",
  1556 => x"862dbdd4",
  1557 => x"08802e88",
  1558 => x"38bdd408",
  1559 => x"519ef72d",
  1560 => x"800bbdd0",
  1561 => x"0cae852d",
  1562 => x"90ae2d02",
  1563 => x"84050d04",
  1564 => x"02fc050d",
  1565 => x"725170fd",
  1566 => x"2ead3870",
  1567 => x"fd248a38",
  1568 => x"70fc2e80",
  1569 => x"c438b1d1",
  1570 => x"0470fe2e",
  1571 => x"b13870ff",
  1572 => x"2e098106",
  1573 => x"bc38bdd0",
  1574 => x"08517080",
  1575 => x"2eb338ff",
  1576 => x"11bdd00c",
  1577 => x"b1d104bd",
  1578 => x"d008f005",
  1579 => x"70bdd00c",
  1580 => x"51708025",
  1581 => x"9c38800b",
  1582 => x"bdd00cb1",
  1583 => x"d104bdd0",
  1584 => x"088105bd",
  1585 => x"d00cb1d1",
  1586 => x"04bdd008",
  1587 => x"9005bdd0",
  1588 => x"0cae852d",
  1589 => x"90ae2d02",
  1590 => x"84050d04",
  1591 => x"02fc050d",
  1592 => x"800bbdd0",
  1593 => x"0cae852d",
  1594 => x"8fc52dbd",
  1595 => x"d408bdc0",
  1596 => x"0cbc9c51",
  1597 => x"91c92d02",
  1598 => x"84050d04",
  1599 => x"7180c4f8",
  1600 => x"0c040000",
  1601 => x"00ffffff",
  1602 => x"ff00ffff",
  1603 => x"ffff00ff",
  1604 => x"ffffff00",
  1605 => x"52657365",
  1606 => x"74000000",
  1607 => x"43617267",
  1608 => x"61722044",
  1609 => x"6973636f",
  1610 => x"2f43696e",
  1611 => x"74612010",
  1612 => x"00000000",
  1613 => x"45786974",
  1614 => x"00000000",
  1615 => x"46444320",
  1616 => x"4f726967",
  1617 => x"696e616c",
  1618 => x"00000000",
  1619 => x"46444320",
  1620 => x"46617374",
  1621 => x"00000000",
  1622 => x"4d756c74",
  1623 => x"69666163",
  1624 => x"65203220",
  1625 => x"456e6162",
  1626 => x"6c656400",
  1627 => x"4d756c74",
  1628 => x"69666163",
  1629 => x"65203220",
  1630 => x"48696464",
  1631 => x"656e0000",
  1632 => x"4d756c74",
  1633 => x"69666163",
  1634 => x"65203220",
  1635 => x"44697361",
  1636 => x"626c6564",
  1637 => x"00000000",
  1638 => x"4d6f7573",
  1639 => x"65204469",
  1640 => x"7361626c",
  1641 => x"65640000",
  1642 => x"4d6f7573",
  1643 => x"6520456e",
  1644 => x"61626c65",
  1645 => x"64000000",
  1646 => x"506c6179",
  1647 => x"63697479",
  1648 => x"20446973",
  1649 => x"61626c65",
  1650 => x"64000000",
  1651 => x"506c6179",
  1652 => x"63697479",
  1653 => x"20456e61",
  1654 => x"626c6564",
  1655 => x"00000000",
  1656 => x"52696768",
  1657 => x"74205368",
  1658 => x"69667420",
  1659 => x"61732042",
  1660 => x"61636b73",
  1661 => x"6c617368",
  1662 => x"00000000",
  1663 => x"52696768",
  1664 => x"74205368",
  1665 => x"69667420",
  1666 => x"61732053",
  1667 => x"68696674",
  1668 => x"00000000",
  1669 => x"536f756e",
  1670 => x"64206f75",
  1671 => x"74707574",
  1672 => x"20537465",
  1673 => x"72656f00",
  1674 => x"536f756e",
  1675 => x"64206f75",
  1676 => x"74707574",
  1677 => x"204d6f6e",
  1678 => x"6f000000",
  1679 => x"54617065",
  1680 => x"20736f75",
  1681 => x"6e642044",
  1682 => x"69736162",
  1683 => x"6c656400",
  1684 => x"54617065",
  1685 => x"20736f75",
  1686 => x"6e642045",
  1687 => x"6e61626c",
  1688 => x"65640000",
  1689 => x"43505520",
  1690 => x"74696d69",
  1691 => x"6e677320",
  1692 => x"4f726967",
  1693 => x"696e616c",
  1694 => x"00000000",
  1695 => x"43505520",
  1696 => x"74696d69",
  1697 => x"6e677320",
  1698 => x"46617374",
  1699 => x"00000000",
  1700 => x"53696e63",
  1701 => x"20736967",
  1702 => x"6e616c73",
  1703 => x"204f7269",
  1704 => x"67696e61",
  1705 => x"6c000000",
  1706 => x"53696e63",
  1707 => x"20736967",
  1708 => x"6e616c73",
  1709 => x"2046696c",
  1710 => x"74657265",
  1711 => x"64000000",
  1712 => x"43525443",
  1713 => x"20547970",
  1714 => x"65203100",
  1715 => x"43525443",
  1716 => x"20547970",
  1717 => x"65203200",
  1718 => x"44697370",
  1719 => x"6c617920",
  1720 => x"436f6c6f",
  1721 => x"72284741",
  1722 => x"29000000",
  1723 => x"44697370",
  1724 => x"6c617920",
  1725 => x"436f6c6f",
  1726 => x"72202841",
  1727 => x"53494329",
  1728 => x"00000000",
  1729 => x"44697370",
  1730 => x"6c617920",
  1731 => x"47726565",
  1732 => x"6e000000",
  1733 => x"44697370",
  1734 => x"6c617920",
  1735 => x"416d6265",
  1736 => x"72000000",
  1737 => x"44697370",
  1738 => x"6c617920",
  1739 => x"4379616e",
  1740 => x"00000000",
  1741 => x"44697370",
  1742 => x"6c617920",
  1743 => x"57686974",
  1744 => x"65000000",
  1745 => x"5363616e",
  1746 => x"6c696e65",
  1747 => x"73204e6f",
  1748 => x"6e650000",
  1749 => x"5363616e",
  1750 => x"6c696e65",
  1751 => x"73204352",
  1752 => x"54203235",
  1753 => x"25000000",
  1754 => x"5363616e",
  1755 => x"6c696e65",
  1756 => x"73204352",
  1757 => x"54203530",
  1758 => x"25000000",
  1759 => x"5363616e",
  1760 => x"6c696e65",
  1761 => x"73204352",
  1762 => x"54203735",
  1763 => x"25000000",
  1764 => x"43617267",
  1765 => x"61204661",
  1766 => x"6c6c6964",
  1767 => x"61000000",
  1768 => x"4f4b0000",
  1769 => x"414d5354",
  1770 => x"52414420",
  1771 => x"44415400",
  1772 => x"16200000",
  1773 => x"14200000",
  1774 => x"15200000",
  1775 => x"53442069",
  1776 => x"6e69742e",
  1777 => x"2e2e0a00",
  1778 => x"53442063",
  1779 => x"61726420",
  1780 => x"72657365",
  1781 => x"74206661",
  1782 => x"696c6564",
  1783 => x"210a0000",
  1784 => x"53444843",
  1785 => x"20657272",
  1786 => x"6f72210a",
  1787 => x"00000000",
  1788 => x"57726974",
  1789 => x"65206661",
  1790 => x"696c6564",
  1791 => x"0a000000",
  1792 => x"52656164",
  1793 => x"20666169",
  1794 => x"6c65640a",
  1795 => x"00000000",
  1796 => x"43617264",
  1797 => x"20696e69",
  1798 => x"74206661",
  1799 => x"696c6564",
  1800 => x"0a000000",
  1801 => x"46415431",
  1802 => x"36202020",
  1803 => x"00000000",
  1804 => x"46415433",
  1805 => x"32202020",
  1806 => x"00000000",
  1807 => x"4e6f2070",
  1808 => x"61727469",
  1809 => x"74696f6e",
  1810 => x"20736967",
  1811 => x"0a000000",
  1812 => x"42616420",
  1813 => x"70617274",
  1814 => x"0a000000",
  1815 => x"4261636b",
  1816 => x"00000000",
  1817 => x"00000002",
  1818 => x"00000002",
  1819 => x"00001914",
  1820 => x"0000034e",
  1821 => x"00000003",
  1822 => x"00001d94",
  1823 => x"00000004",
  1824 => x"00000003",
  1825 => x"00001d7c",
  1826 => x"00000006",
  1827 => x"00000003",
  1828 => x"00001d74",
  1829 => x"00000002",
  1830 => x"00000003",
  1831 => x"00001d6c",
  1832 => x"00000002",
  1833 => x"00000003",
  1834 => x"00001d64",
  1835 => x"00000002",
  1836 => x"00000003",
  1837 => x"00001d5c",
  1838 => x"00000002",
  1839 => x"00000003",
  1840 => x"00001d54",
  1841 => x"00000002",
  1842 => x"00000003",
  1843 => x"00001d4c",
  1844 => x"00000002",
  1845 => x"00000003",
  1846 => x"00001d44",
  1847 => x"00000002",
  1848 => x"00000003",
  1849 => x"00001d3c",
  1850 => x"00000002",
  1851 => x"00000003",
  1852 => x"00001d30",
  1853 => x"00000003",
  1854 => x"00000003",
  1855 => x"00001d28",
  1856 => x"00000002",
  1857 => x"00000002",
  1858 => x"0000191c",
  1859 => x"000018dc",
  1860 => x"00000002",
  1861 => x"00001934",
  1862 => x"000007cc",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"00000000",
  1866 => x"0000193c",
  1867 => x"0000194c",
  1868 => x"00001958",
  1869 => x"0000196c",
  1870 => x"00001980",
  1871 => x"00001998",
  1872 => x"000019a8",
  1873 => x"000019b8",
  1874 => x"000019cc",
  1875 => x"000019e0",
  1876 => x"000019fc",
  1877 => x"00001a14",
  1878 => x"00001a28",
  1879 => x"00001a3c",
  1880 => x"00001a50",
  1881 => x"00001a64",
  1882 => x"00001a7c",
  1883 => x"00001a90",
  1884 => x"00001aa8",
  1885 => x"00001ac0",
  1886 => x"00001acc",
  1887 => x"00001ad8",
  1888 => x"00001aec",
  1889 => x"00001b04",
  1890 => x"00001b14",
  1891 => x"00001b24",
  1892 => x"00001b34",
  1893 => x"00001b44",
  1894 => x"00001b54",
  1895 => x"00001b68",
  1896 => x"00001b7c",
  1897 => x"00000004",
  1898 => x"00001b90",
  1899 => x"00001da4",
  1900 => x"00000004",
  1901 => x"00001ba0",
  1902 => x"00001c68",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000000",
  1913 => x"00000000",
  1914 => x"00000000",
  1915 => x"00000000",
  1916 => x"00000000",
  1917 => x"00000000",
  1918 => x"00000000",
  1919 => x"00000000",
  1920 => x"00000000",
  1921 => x"00000000",
  1922 => x"00000000",
  1923 => x"00000000",
  1924 => x"00000000",
  1925 => x"00000000",
  1926 => x"00000000",
  1927 => x"00000002",
  1928 => x"0000227c",
  1929 => x"000016d0",
  1930 => x"00000002",
  1931 => x"0000229a",
  1932 => x"000016d0",
  1933 => x"00000002",
  1934 => x"000022b8",
  1935 => x"000016d0",
  1936 => x"00000002",
  1937 => x"000022d6",
  1938 => x"000016d0",
  1939 => x"00000002",
  1940 => x"000022f4",
  1941 => x"000016d0",
  1942 => x"00000002",
  1943 => x"00002312",
  1944 => x"000016d0",
  1945 => x"00000002",
  1946 => x"00002330",
  1947 => x"000016d0",
  1948 => x"00000002",
  1949 => x"0000234e",
  1950 => x"000016d0",
  1951 => x"00000002",
  1952 => x"0000236c",
  1953 => x"000016d0",
  1954 => x"00000002",
  1955 => x"0000238a",
  1956 => x"000016d0",
  1957 => x"00000002",
  1958 => x"000023a8",
  1959 => x"000016d0",
  1960 => x"00000002",
  1961 => x"000023c6",
  1962 => x"000016d0",
  1963 => x"00000002",
  1964 => x"000023e4",
  1965 => x"000016d0",
  1966 => x"00000004",
  1967 => x"00001c5c",
  1968 => x"00000000",
  1969 => x"00000000",
  1970 => x"00000000",
  1971 => x"00001870",
  1972 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

