-- ZPU
--
-- Copyright 2004-2008 oharboe - �yvind Harboe - oyvind.harboe@zylin.com
-- Modified by Alastair M. Robinson for the ZPUFlex project.
--
-- The FreeBSD license
-- 
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimer in the documentation and/or other materials
--    provided with the distribution.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE ZPU PROJECT ``AS IS'' AND ANY
-- EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO,
-- THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A
-- PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE
-- ZPU PROJECT OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT,
-- INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT,
-- STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE)
-- ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF
-- ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
-- 
-- The views and conclusions contained in the software and documentation
-- are those of the authors and should not be interpreted as representing
-- official policies, either expressed or implied, of the ZPU Project.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;

entity CtrlROM_ROM is
generic
	(
		maxAddrBitBRAM : integer := maxAddrBitBRAMLimit -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	areset : in std_logic := '0';
	from_zpu : in ZPU_ToROM;
	to_zpu : out ZPU_FromROM
);
end CtrlROM_ROM;

architecture arch of CtrlROM_ROM is

type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(wordSize-1 downto 0);

shared variable ram : ram_type :=
(
     0 => x"0b0b0b0b",
     1 => x"8c0b0b0b",
     2 => x"0b81e004",
     3 => x"0b0b0b0b",
     4 => x"8c04ff0d",
     5 => x"80040400",
     6 => x"00000016",
     7 => x"00000000",
     8 => x"0b0b0bbd",
     9 => x"98080b0b",
    10 => x"0bbd9c08",
    11 => x"0b0b0bbd",
    12 => x"a0080b0b",
    13 => x"0b0b9808",
    14 => x"2d0b0b0b",
    15 => x"bda00c0b",
    16 => x"0b0bbd9c",
    17 => x"0c0b0b0b",
    18 => x"bd980c04",
    19 => x"00000000",
    20 => x"00000000",
    21 => x"00000000",
    22 => x"00000000",
    23 => x"00000000",
    24 => x"71fd0608",
    25 => x"72830609",
    26 => x"81058205",
    27 => x"832b2a83",
    28 => x"ffff0652",
    29 => x"0471fc06",
    30 => x"08728306",
    31 => x"09810583",
    32 => x"05101010",
    33 => x"2a81ff06",
    34 => x"520471fd",
    35 => x"060883ff",
    36 => x"ff738306",
    37 => x"09810582",
    38 => x"05832b2b",
    39 => x"09067383",
    40 => x"ffff0673",
    41 => x"83060981",
    42 => x"05820583",
    43 => x"2b0b2b07",
    44 => x"72fc060c",
    45 => x"51510471",
    46 => x"fc06080b",
    47 => x"0b0bb1c8",
    48 => x"73830610",
    49 => x"10050806",
    50 => x"7381ff06",
    51 => x"73830609",
    52 => x"81058305",
    53 => x"1010102b",
    54 => x"0772fc06",
    55 => x"0c515104",
    56 => x"bd987080",
    57 => x"c7c8278b",
    58 => x"38807170",
    59 => x"8405530c",
    60 => x"81e2048c",
    61 => x"5188c504",
    62 => x"02fc050d",
    63 => x"f880518f",
    64 => x"0bbda80c",
    65 => x"9f0bbdac",
    66 => x"0ca07170",
    67 => x"81055334",
    68 => x"bdac08ff",
    69 => x"05bdac0c",
    70 => x"bdac0880",
    71 => x"25eb38bd",
    72 => x"a808ff05",
    73 => x"bda80cbd",
    74 => x"a8088025",
    75 => x"d738800b",
    76 => x"bdac0c80",
    77 => x"0bbda80c",
    78 => x"0284050d",
    79 => x"0402f005",
    80 => x"0df88053",
    81 => x"f8a05483",
    82 => x"bf527370",
    83 => x"81055533",
    84 => x"51707370",
    85 => x"81055534",
    86 => x"ff125271",
    87 => x"8025eb38",
    88 => x"fbc0539f",
    89 => x"52a07370",
    90 => x"81055534",
    91 => x"ff125271",
    92 => x"8025f238",
    93 => x"0290050d",
    94 => x"0402f405",
    95 => x"0d74538e",
    96 => x"0bbda808",
    97 => x"258f3882",
    98 => x"bd2dbda8",
    99 => x"08ff05bd",
   100 => x"a80c82ff",
   101 => x"04bda808",
   102 => x"bdac0853",
   103 => x"51728a2e",
   104 => x"098106b7",
   105 => x"38715171",
   106 => x"9f24a038",
   107 => x"bda808a0",
   108 => x"2911f880",
   109 => x"115151a0",
   110 => x"7134bdac",
   111 => x"088105bd",
   112 => x"ac0cbdac",
   113 => x"08519f71",
   114 => x"25e23880",
   115 => x"0bbdac0c",
   116 => x"bda80881",
   117 => x"05bda80c",
   118 => x"83ef0470",
   119 => x"a02912f8",
   120 => x"80115151",
   121 => x"727134bd",
   122 => x"ac088105",
   123 => x"bdac0cbd",
   124 => x"ac08a02e",
   125 => x"0981068e",
   126 => x"38800bbd",
   127 => x"ac0cbda8",
   128 => x"088105bd",
   129 => x"a80c028c",
   130 => x"050d0402",
   131 => x"e8050d77",
   132 => x"79565688",
   133 => x"0bfc1677",
   134 => x"712c8f06",
   135 => x"54525480",
   136 => x"53727225",
   137 => x"95387153",
   138 => x"fbe01451",
   139 => x"87713481",
   140 => x"14ff1454",
   141 => x"5472f138",
   142 => x"7153f915",
   143 => x"76712c87",
   144 => x"06535171",
   145 => x"802e8b38",
   146 => x"fbe01451",
   147 => x"71713481",
   148 => x"1454728e",
   149 => x"2495388f",
   150 => x"733153fb",
   151 => x"e01451a0",
   152 => x"71348114",
   153 => x"ff145454",
   154 => x"72f13802",
   155 => x"98050d04",
   156 => x"02ec050d",
   157 => x"800bbdb0",
   158 => x"0cf68c08",
   159 => x"f6900871",
   160 => x"882c5654",
   161 => x"81ff0652",
   162 => x"73722588",
   163 => x"38715482",
   164 => x"0bbdb00c",
   165 => x"72882c73",
   166 => x"81ff0654",
   167 => x"55747325",
   168 => x"8b3872bd",
   169 => x"b0088407",
   170 => x"bdb00c55",
   171 => x"73842b86",
   172 => x"a0712583",
   173 => x"7131700b",
   174 => x"0b0bb8a8",
   175 => x"0c81712b",
   176 => x"ff05f688",
   177 => x"0cfdfc13",
   178 => x"ff122c78",
   179 => x"8829ff94",
   180 => x"0570812c",
   181 => x"bdb00852",
   182 => x"58525551",
   183 => x"52547680",
   184 => x"2e853870",
   185 => x"81075170",
   186 => x"f6940c71",
   187 => x"098105f6",
   188 => x"800c7209",
   189 => x"8105f684",
   190 => x"0c029405",
   191 => x"0d0402f4",
   192 => x"050d7453",
   193 => x"72708105",
   194 => x"5480f52d",
   195 => x"5271802e",
   196 => x"89387151",
   197 => x"82f92d86",
   198 => x"8404810b",
   199 => x"bd980c02",
   200 => x"8c050d04",
   201 => x"02fc050d",
   202 => x"81808051",
   203 => x"c0115170",
   204 => x"fb380284",
   205 => x"050d0402",
   206 => x"fc050d84",
   207 => x"bf5186a4",
   208 => x"2dff1151",
   209 => x"708025f6",
   210 => x"38028405",
   211 => x"0d0402fc",
   212 => x"050dec51",
   213 => x"83710c86",
   214 => x"a42d8271",
   215 => x"0c028405",
   216 => x"0d0402fc",
   217 => x"050dec51",
   218 => x"92710c86",
   219 => x"a42d8271",
   220 => x"0c028405",
   221 => x"0d0402dc",
   222 => x"050d7a54",
   223 => x"807453bd",
   224 => x"b45259a8",
   225 => x"e72dbd98",
   226 => x"08792e81",
   227 => x"9138bdb8",
   228 => x"0870f80c",
   229 => x"891580f5",
   230 => x"2d8a1680",
   231 => x"f52d7182",
   232 => x"80290588",
   233 => x"1780f52d",
   234 => x"70848080",
   235 => x"2912f40c",
   236 => x"57555755",
   237 => x"a40bec0c",
   238 => x"78ff1655",
   239 => x"5873792e",
   240 => x"8b388118",
   241 => x"74812a55",
   242 => x"5873f738",
   243 => x"f7185881",
   244 => x"59807525",
   245 => x"80c83877",
   246 => x"52735184",
   247 => x"8b2dbe80",
   248 => x"52bdb451",
   249 => x"aba62dbd",
   250 => x"9808802e",
   251 => x"9a38be80",
   252 => x"5783fc56",
   253 => x"76708405",
   254 => x"5808e80c",
   255 => x"fc165675",
   256 => x"8025f138",
   257 => x"888e04bd",
   258 => x"98085984",
   259 => x"8055bdb4",
   260 => x"51aaf82d",
   261 => x"fc801581",
   262 => x"15555587",
   263 => x"d10486b7",
   264 => x"2d840bec",
   265 => x"0c78802e",
   266 => x"8d38b8ac",
   267 => x"51918d2d",
   268 => x"8f902d88",
   269 => x"bc04bae8",
   270 => x"51918d2d",
   271 => x"78bd980c",
   272 => x"02a4050d",
   273 => x"0402e005",
   274 => x"0d805584",
   275 => x"0bec0c8e",
   276 => x"f12d8bdb",
   277 => x"2d81f82d",
   278 => x"9fdc2dbd",
   279 => x"9808752e",
   280 => x"82e4388c",
   281 => x"0bec0cb6",
   282 => x"e852bdb4",
   283 => x"51a8e72d",
   284 => x"bd980875",
   285 => x"2e80e538",
   286 => x"bdb80875",
   287 => x"ff125659",
   288 => x"5673752e",
   289 => x"8b388118",
   290 => x"74812a55",
   291 => x"5873f738",
   292 => x"f7185880",
   293 => x"762580c4",
   294 => x"38775273",
   295 => x"51848b2d",
   296 => x"be8052bd",
   297 => x"b451aba6",
   298 => x"2dbd9808",
   299 => x"802e9a38",
   300 => x"be805783",
   301 => x"fc557670",
   302 => x"84055808",
   303 => x"e80cfc15",
   304 => x"55748025",
   305 => x"f13889cc",
   306 => x"04848056",
   307 => x"bdb451aa",
   308 => x"f82dfc80",
   309 => x"16811555",
   310 => x"56899304",
   311 => x"bdb808f8",
   312 => x"0c86b72d",
   313 => x"840bec0c",
   314 => x"86f651b1",
   315 => x"c02db8ac",
   316 => x"51918d2d",
   317 => x"8f902d8b",
   318 => x"e72d919d",
   319 => x"2db8cc0b",
   320 => x"80f52d70",
   321 => x"822b9c06",
   322 => x"b8c00b80",
   323 => x"f52d8306",
   324 => x"7107b8d8",
   325 => x"0b80f52d",
   326 => x"70852ba0",
   327 => x"06b8e40b",
   328 => x"80f52d70",
   329 => x"862b80c0",
   330 => x"06747307",
   331 => x"07b8f00b",
   332 => x"80f52d70",
   333 => x"872b8180",
   334 => x"06b8fc0b",
   335 => x"80f52d70",
   336 => x"882b8280",
   337 => x"06747307",
   338 => x"07b9880b",
   339 => x"80f52d70",
   340 => x"892b8480",
   341 => x"06b9940b",
   342 => x"80f52d70",
   343 => x"8a2b8880",
   344 => x"06747307",
   345 => x"07b9a00b",
   346 => x"80f52d70",
   347 => x"8b2b9080",
   348 => x"06b9ac0b",
   349 => x"80f52d70",
   350 => x"8c2ba080",
   351 => x"06747307",
   352 => x"07b9b80b",
   353 => x"80f52d70",
   354 => x"8d2b81c0",
   355 => x"8006b9c4",
   356 => x"0b80f52d",
   357 => x"708f2b82",
   358 => x"80800674",
   359 => x"730707fc",
   360 => x"0c545454",
   361 => x"54545454",
   362 => x"54545454",
   363 => x"54545454",
   364 => x"545b5452",
   365 => x"57545486",
   366 => x"53bd9808",
   367 => x"83388453",
   368 => x"72ec0c89",
   369 => x"f704800b",
   370 => x"bd980c02",
   371 => x"a0050d04",
   372 => x"71980c04",
   373 => x"ffb008bd",
   374 => x"980c0481",
   375 => x"0bffb00c",
   376 => x"04800bff",
   377 => x"b00c0402",
   378 => x"f4050d8c",
   379 => x"e904bd98",
   380 => x"0881f02e",
   381 => x"09810689",
   382 => x"38810bbb",
   383 => x"cc0c8ce9",
   384 => x"04bd9808",
   385 => x"81e02e09",
   386 => x"81068938",
   387 => x"810bbbd0",
   388 => x"0c8ce904",
   389 => x"bd980852",
   390 => x"bbd00880",
   391 => x"2e8838bd",
   392 => x"98088180",
   393 => x"05527184",
   394 => x"2c728f06",
   395 => x"5353bbcc",
   396 => x"08802e99",
   397 => x"38728429",
   398 => x"bb8c0572",
   399 => x"1381712b",
   400 => x"70097308",
   401 => x"06730c51",
   402 => x"53538cdf",
   403 => x"04728429",
   404 => x"bb8c0572",
   405 => x"1383712b",
   406 => x"72080772",
   407 => x"0c535380",
   408 => x"0bbbd00c",
   409 => x"800bbbcc",
   410 => x"0cbdc051",
   411 => x"8dea2dbd",
   412 => x"9808ff24",
   413 => x"fef83880",
   414 => x"0bbd980c",
   415 => x"028c050d",
   416 => x"0402f805",
   417 => x"0dbb8c52",
   418 => x"8f518072",
   419 => x"70840554",
   420 => x"0cff1151",
   421 => x"708025f2",
   422 => x"38028805",
   423 => x"0d0402f0",
   424 => x"050d7551",
   425 => x"8be12d70",
   426 => x"822cfc06",
   427 => x"bb8c1172",
   428 => x"109e0671",
   429 => x"0870722a",
   430 => x"70830682",
   431 => x"742b7009",
   432 => x"7406760c",
   433 => x"54515657",
   434 => x"5351538b",
   435 => x"db2d71bd",
   436 => x"980c0290",
   437 => x"050d0402",
   438 => x"fc050d72",
   439 => x"5180710c",
   440 => x"800b8412",
   441 => x"0c028405",
   442 => x"0d0402f0",
   443 => x"050d7570",
   444 => x"08841208",
   445 => x"535353ff",
   446 => x"5471712e",
   447 => x"a8388be1",
   448 => x"2d841308",
   449 => x"70842914",
   450 => x"88117008",
   451 => x"7081ff06",
   452 => x"84180881",
   453 => x"11870684",
   454 => x"1a0c5351",
   455 => x"55515151",
   456 => x"8bdb2d71",
   457 => x"5473bd98",
   458 => x"0c029005",
   459 => x"0d0402f8",
   460 => x"050d8be1",
   461 => x"2de00870",
   462 => x"8b2a7081",
   463 => x"06515252",
   464 => x"70802e9d",
   465 => x"38bdc008",
   466 => x"708429bd",
   467 => x"c8057381",
   468 => x"ff06710c",
   469 => x"5151bdc0",
   470 => x"08811187",
   471 => x"06bdc00c",
   472 => x"51800bbd",
   473 => x"e80c8bd4",
   474 => x"2d8bdb2d",
   475 => x"0288050d",
   476 => x"0402fc05",
   477 => x"0dbdc051",
   478 => x"8dd72d8d",
   479 => x"812d8eae",
   480 => x"518bd02d",
   481 => x"0284050d",
   482 => x"04bdec08",
   483 => x"bd980c04",
   484 => x"02fc050d",
   485 => x"8f9a048b",
   486 => x"e72d80f6",
   487 => x"518d9e2d",
   488 => x"bd9808f3",
   489 => x"3880da51",
   490 => x"8d9e2dbd",
   491 => x"9808e838",
   492 => x"bd9808bb",
   493 => x"d80cbd98",
   494 => x"085184f0",
   495 => x"2d028405",
   496 => x"0d0402ec",
   497 => x"050d7654",
   498 => x"8052870b",
   499 => x"881580f5",
   500 => x"2d565374",
   501 => x"72248338",
   502 => x"a0537251",
   503 => x"82f92d81",
   504 => x"128b1580",
   505 => x"f52d5452",
   506 => x"727225de",
   507 => x"38029405",
   508 => x"0d0402f0",
   509 => x"050dbdec",
   510 => x"085481f8",
   511 => x"2d800bbd",
   512 => x"f00c7308",
   513 => x"802e8180",
   514 => x"38820bbd",
   515 => x"ac0cbdf0",
   516 => x"088f06bd",
   517 => x"a80c7308",
   518 => x"5271832e",
   519 => x"96387183",
   520 => x"26893871",
   521 => x"812eaf38",
   522 => x"90f30471",
   523 => x"852e9f38",
   524 => x"90f30488",
   525 => x"1480f52d",
   526 => x"841508b6",
   527 => x"f4535452",
   528 => x"85fe2d71",
   529 => x"84291370",
   530 => x"08525290",
   531 => x"f7047351",
   532 => x"8fc22d90",
   533 => x"f304bbd4",
   534 => x"08881508",
   535 => x"2c708106",
   536 => x"51527180",
   537 => x"2e8738b6",
   538 => x"f85190f0",
   539 => x"04b6fc51",
   540 => x"85fe2d84",
   541 => x"14085185",
   542 => x"fe2dbdf0",
   543 => x"088105bd",
   544 => x"f00c8c14",
   545 => x"54908204",
   546 => x"0290050d",
   547 => x"0471bdec",
   548 => x"0c8ff22d",
   549 => x"bdf008ff",
   550 => x"05bdf40c",
   551 => x"0402e805",
   552 => x"0dbdec08",
   553 => x"bdf80857",
   554 => x"5587518d",
   555 => x"9e2dbd98",
   556 => x"08812a70",
   557 => x"81065152",
   558 => x"71802ea0",
   559 => x"3891c304",
   560 => x"8be72d87",
   561 => x"518d9e2d",
   562 => x"bd9808f4",
   563 => x"38bbd808",
   564 => x"813270bb",
   565 => x"d80c7052",
   566 => x"5284f02d",
   567 => x"80fe518d",
   568 => x"9e2dbd98",
   569 => x"08802ea6",
   570 => x"38bbd808",
   571 => x"802e9138",
   572 => x"800bbbd8",
   573 => x"0c805184",
   574 => x"f02d9280",
   575 => x"048be72d",
   576 => x"80fe518d",
   577 => x"9e2dbd98",
   578 => x"08f33886",
   579 => x"e22dbbd8",
   580 => x"08903881",
   581 => x"fd518d9e",
   582 => x"2d81fa51",
   583 => x"8d9e2d97",
   584 => x"d30481f5",
   585 => x"518d9e2d",
   586 => x"bd980881",
   587 => x"2a708106",
   588 => x"51527180",
   589 => x"2eaf38bd",
   590 => x"f4085271",
   591 => x"802e8938",
   592 => x"ff12bdf4",
   593 => x"0c92e504",
   594 => x"bdf00810",
   595 => x"bdf00805",
   596 => x"70842916",
   597 => x"51528812",
   598 => x"08802e89",
   599 => x"38ff5188",
   600 => x"12085271",
   601 => x"2d81f251",
   602 => x"8d9e2dbd",
   603 => x"9808812a",
   604 => x"70810651",
   605 => x"5271802e",
   606 => x"b138bdf0",
   607 => x"08ff11bd",
   608 => x"f4085653",
   609 => x"53737225",
   610 => x"89388114",
   611 => x"bdf40c93",
   612 => x"aa047210",
   613 => x"13708429",
   614 => x"16515288",
   615 => x"1208802e",
   616 => x"8938fe51",
   617 => x"88120852",
   618 => x"712d81fd",
   619 => x"518d9e2d",
   620 => x"bd980881",
   621 => x"2a708106",
   622 => x"51527180",
   623 => x"2ead38bd",
   624 => x"f408802e",
   625 => x"8938800b",
   626 => x"bdf40c93",
   627 => x"eb04bdf0",
   628 => x"0810bdf0",
   629 => x"08057084",
   630 => x"29165152",
   631 => x"88120880",
   632 => x"2e8938fd",
   633 => x"51881208",
   634 => x"52712d81",
   635 => x"fa518d9e",
   636 => x"2dbd9808",
   637 => x"812a7081",
   638 => x"06515271",
   639 => x"802eae38",
   640 => x"bdf008ff",
   641 => x"115452bd",
   642 => x"f4087325",
   643 => x"883872bd",
   644 => x"f40c94ad",
   645 => x"04711012",
   646 => x"70842916",
   647 => x"51528812",
   648 => x"08802e89",
   649 => x"38fc5188",
   650 => x"12085271",
   651 => x"2dbdf408",
   652 => x"70535473",
   653 => x"802e8a38",
   654 => x"8c15ff15",
   655 => x"555594b3",
   656 => x"04820bbd",
   657 => x"ac0c718f",
   658 => x"06bda80c",
   659 => x"81eb518d",
   660 => x"9e2dbd98",
   661 => x"08812a70",
   662 => x"81065152",
   663 => x"71802ead",
   664 => x"38740885",
   665 => x"2e098106",
   666 => x"a4388815",
   667 => x"80f52dff",
   668 => x"05527188",
   669 => x"1681b72d",
   670 => x"71982b52",
   671 => x"71802588",
   672 => x"38800b88",
   673 => x"1681b72d",
   674 => x"74518fc2",
   675 => x"2d81f451",
   676 => x"8d9e2dbd",
   677 => x"9808812a",
   678 => x"70810651",
   679 => x"5271802e",
   680 => x"b3387408",
   681 => x"852e0981",
   682 => x"06aa3888",
   683 => x"1580f52d",
   684 => x"81055271",
   685 => x"881681b7",
   686 => x"2d7181ff",
   687 => x"068b1680",
   688 => x"f52d5452",
   689 => x"72722787",
   690 => x"38728816",
   691 => x"81b72d74",
   692 => x"518fc22d",
   693 => x"80da518d",
   694 => x"9e2dbd98",
   695 => x"08812a70",
   696 => x"81065152",
   697 => x"71802e81",
   698 => x"a638bdec",
   699 => x"08bdf408",
   700 => x"55537380",
   701 => x"2e8a388c",
   702 => x"13ff1555",
   703 => x"5395f204",
   704 => x"72085271",
   705 => x"822ea638",
   706 => x"71822689",
   707 => x"3871812e",
   708 => x"a938978f",
   709 => x"0471832e",
   710 => x"b1387184",
   711 => x"2e098106",
   712 => x"80ed3888",
   713 => x"13085191",
   714 => x"8d2d978f",
   715 => x"04bdf408",
   716 => x"51881308",
   717 => x"52712d97",
   718 => x"8f04810b",
   719 => x"8814082b",
   720 => x"bbd40832",
   721 => x"bbd40c96",
   722 => x"e5048813",
   723 => x"80f52d81",
   724 => x"058b1480",
   725 => x"f52d5354",
   726 => x"71742483",
   727 => x"38805473",
   728 => x"881481b7",
   729 => x"2d8ff22d",
   730 => x"978f0475",
   731 => x"08802ea2",
   732 => x"38750851",
   733 => x"8d9e2dbd",
   734 => x"98088106",
   735 => x"5271802e",
   736 => x"8b38bdf4",
   737 => x"08518416",
   738 => x"0852712d",
   739 => x"88165675",
   740 => x"da388054",
   741 => x"800bbdac",
   742 => x"0c738f06",
   743 => x"bda80ca0",
   744 => x"5273bdf4",
   745 => x"082e0981",
   746 => x"069838bd",
   747 => x"f008ff05",
   748 => x"74327009",
   749 => x"81057072",
   750 => x"079f2a91",
   751 => x"71315151",
   752 => x"53537151",
   753 => x"82f92d81",
   754 => x"14548e74",
   755 => x"25c638bb",
   756 => x"d8085271",
   757 => x"bd980c02",
   758 => x"98050d04",
   759 => x"02f4050d",
   760 => x"d45281ff",
   761 => x"720c7108",
   762 => x"5381ff72",
   763 => x"0c72882b",
   764 => x"83fe8006",
   765 => x"72087081",
   766 => x"ff065152",
   767 => x"5381ff72",
   768 => x"0c727107",
   769 => x"882b7208",
   770 => x"7081ff06",
   771 => x"51525381",
   772 => x"ff720c72",
   773 => x"7107882b",
   774 => x"72087081",
   775 => x"ff067207",
   776 => x"bd980c52",
   777 => x"53028c05",
   778 => x"0d0402f4",
   779 => x"050d7476",
   780 => x"7181ff06",
   781 => x"d40c5353",
   782 => x"bdfc0885",
   783 => x"3871892b",
   784 => x"5271982a",
   785 => x"d40c7190",
   786 => x"2a7081ff",
   787 => x"06d40c51",
   788 => x"71882a70",
   789 => x"81ff06d4",
   790 => x"0c517181",
   791 => x"ff06d40c",
   792 => x"72902a70",
   793 => x"81ff06d4",
   794 => x"0c51d408",
   795 => x"7081ff06",
   796 => x"515182b8",
   797 => x"bf527081",
   798 => x"ff2e0981",
   799 => x"06943881",
   800 => x"ff0bd40c",
   801 => x"d4087081",
   802 => x"ff06ff14",
   803 => x"54515171",
   804 => x"e53870bd",
   805 => x"980c028c",
   806 => x"050d0402",
   807 => x"fc050d81",
   808 => x"c75181ff",
   809 => x"0bd40cff",
   810 => x"11517080",
   811 => x"25f43802",
   812 => x"84050d04",
   813 => x"02f4050d",
   814 => x"81ff0bd4",
   815 => x"0c935380",
   816 => x"5287fc80",
   817 => x"c15198aa",
   818 => x"2dbd9808",
   819 => x"8b3881ff",
   820 => x"0bd40c81",
   821 => x"5399e104",
   822 => x"999b2dff",
   823 => x"135372df",
   824 => x"3872bd98",
   825 => x"0c028c05",
   826 => x"0d0402ec",
   827 => x"050d810b",
   828 => x"bdfc0c84",
   829 => x"54d00870",
   830 => x"8f2a7081",
   831 => x"06515153",
   832 => x"72f33872",
   833 => x"d00c999b",
   834 => x"2db78051",
   835 => x"85fe2dd0",
   836 => x"08708f2a",
   837 => x"70810651",
   838 => x"515372f3",
   839 => x"38810bd0",
   840 => x"0cb15380",
   841 => x"5284d480",
   842 => x"c05198aa",
   843 => x"2dbd9808",
   844 => x"812e9338",
   845 => x"72822ebd",
   846 => x"38ff1353",
   847 => x"72e538ff",
   848 => x"145473ff",
   849 => x"b038999b",
   850 => x"2d83aa52",
   851 => x"849c80c8",
   852 => x"5198aa2d",
   853 => x"bd980881",
   854 => x"2e098106",
   855 => x"923897dc",
   856 => x"2dbd9808",
   857 => x"83ffff06",
   858 => x"537283aa",
   859 => x"2e9d3899",
   860 => x"b42d9b86",
   861 => x"04b78c51",
   862 => x"85fe2d80",
   863 => x"539cd404",
   864 => x"b7a45185",
   865 => x"fe2d8054",
   866 => x"9ca60481",
   867 => x"ff0bd40c",
   868 => x"b154999b",
   869 => x"2d8fcf53",
   870 => x"805287fc",
   871 => x"80f75198",
   872 => x"aa2dbd98",
   873 => x"0855bd98",
   874 => x"08812e09",
   875 => x"81069b38",
   876 => x"81ff0bd4",
   877 => x"0c820a52",
   878 => x"849c80e9",
   879 => x"5198aa2d",
   880 => x"bd980880",
   881 => x"2e8d3899",
   882 => x"9b2dff13",
   883 => x"5372c938",
   884 => x"9c990481",
   885 => x"ff0bd40c",
   886 => x"bd980852",
   887 => x"87fc80fa",
   888 => x"5198aa2d",
   889 => x"bd9808b1",
   890 => x"3881ff0b",
   891 => x"d40cd408",
   892 => x"5381ff0b",
   893 => x"d40c81ff",
   894 => x"0bd40c81",
   895 => x"ff0bd40c",
   896 => x"81ff0bd4",
   897 => x"0c72862a",
   898 => x"70810676",
   899 => x"56515372",
   900 => x"9538bd98",
   901 => x"08549ca6",
   902 => x"0473822e",
   903 => x"fee238ff",
   904 => x"145473fe",
   905 => x"ed3873bd",
   906 => x"fc0c738b",
   907 => x"38815287",
   908 => x"fc80d051",
   909 => x"98aa2d81",
   910 => x"ff0bd40c",
   911 => x"d008708f",
   912 => x"2a708106",
   913 => x"51515372",
   914 => x"f33872d0",
   915 => x"0c81ff0b",
   916 => x"d40c8153",
   917 => x"72bd980c",
   918 => x"0294050d",
   919 => x"0402e805",
   920 => x"0d785580",
   921 => x"5681ff0b",
   922 => x"d40cd008",
   923 => x"708f2a70",
   924 => x"81065151",
   925 => x"5372f338",
   926 => x"82810bd0",
   927 => x"0c81ff0b",
   928 => x"d40c7752",
   929 => x"87fc80d1",
   930 => x"5198aa2d",
   931 => x"80dbc6df",
   932 => x"54bd9808",
   933 => x"802e8a38",
   934 => x"b7c45185",
   935 => x"fe2d9df4",
   936 => x"0481ff0b",
   937 => x"d40cd408",
   938 => x"7081ff06",
   939 => x"51537281",
   940 => x"fe2e0981",
   941 => x"069d3880",
   942 => x"ff5397dc",
   943 => x"2dbd9808",
   944 => x"75708405",
   945 => x"570cff13",
   946 => x"53728025",
   947 => x"ed388156",
   948 => x"9dd904ff",
   949 => x"145473c9",
   950 => x"3881ff0b",
   951 => x"d40c81ff",
   952 => x"0bd40cd0",
   953 => x"08708f2a",
   954 => x"70810651",
   955 => x"515372f3",
   956 => x"3872d00c",
   957 => x"75bd980c",
   958 => x"0298050d",
   959 => x"0402e805",
   960 => x"0d77797b",
   961 => x"58555580",
   962 => x"53727625",
   963 => x"a3387470",
   964 => x"81055680",
   965 => x"f52d7470",
   966 => x"81055680",
   967 => x"f52d5252",
   968 => x"71712e86",
   969 => x"3881519e",
   970 => x"b2048113",
   971 => x"539e8904",
   972 => x"805170bd",
   973 => x"980c0298",
   974 => x"050d0402",
   975 => x"ec050d76",
   976 => x"5574802e",
   977 => x"be389a15",
   978 => x"80e02d51",
   979 => x"abff2dbd",
   980 => x"9808bd98",
   981 => x"0880c4b0",
   982 => x"0cbd9808",
   983 => x"545480c4",
   984 => x"8c08802e",
   985 => x"99389415",
   986 => x"80e02d51",
   987 => x"abff2dbd",
   988 => x"9808902b",
   989 => x"83fff00a",
   990 => x"06707507",
   991 => x"51537280",
   992 => x"c4b00c80",
   993 => x"c4b00853",
   994 => x"72802e9d",
   995 => x"3880c484",
   996 => x"08fe1471",
   997 => x"2980c498",
   998 => x"080580c4",
   999 => x"b40c7084",
  1000 => x"2b80c490",
  1001 => x"0c549fd7",
  1002 => x"0480c49c",
  1003 => x"0880c4b0",
  1004 => x"0c80c4a0",
  1005 => x"0880c4b4",
  1006 => x"0c80c48c",
  1007 => x"08802e8b",
  1008 => x"3880c484",
  1009 => x"08842b53",
  1010 => x"9fd20480",
  1011 => x"c4a40884",
  1012 => x"2b537280",
  1013 => x"c4900c02",
  1014 => x"94050d04",
  1015 => x"02d8050d",
  1016 => x"800b80c4",
  1017 => x"8c0c8454",
  1018 => x"99ea2dbd",
  1019 => x"9808802e",
  1020 => x"9538be80",
  1021 => x"5280519c",
  1022 => x"dd2dbd98",
  1023 => x"08802e86",
  1024 => x"38fe54a0",
  1025 => x"8e04ff14",
  1026 => x"54738024",
  1027 => x"db38738c",
  1028 => x"38b7d451",
  1029 => x"85fe2d73",
  1030 => x"55a5b804",
  1031 => x"8056810b",
  1032 => x"80c4b80c",
  1033 => x"8853b7e8",
  1034 => x"52beb651",
  1035 => x"9dfd2dbd",
  1036 => x"9808762e",
  1037 => x"09810688",
  1038 => x"38bd9808",
  1039 => x"80c4b80c",
  1040 => x"8853b7f4",
  1041 => x"52bed251",
  1042 => x"9dfd2dbd",
  1043 => x"98088838",
  1044 => x"bd980880",
  1045 => x"c4b80c80",
  1046 => x"c4b80880",
  1047 => x"2e80fc38",
  1048 => x"80c1c60b",
  1049 => x"80f52d80",
  1050 => x"c1c70b80",
  1051 => x"f52d7198",
  1052 => x"2b71902b",
  1053 => x"0780c1c8",
  1054 => x"0b80f52d",
  1055 => x"70882b72",
  1056 => x"0780c1c9",
  1057 => x"0b80f52d",
  1058 => x"710780c1",
  1059 => x"fe0b80f5",
  1060 => x"2d80c1ff",
  1061 => x"0b80f52d",
  1062 => x"71882b07",
  1063 => x"535f5452",
  1064 => x"5a565755",
  1065 => x"7381abaa",
  1066 => x"2e098106",
  1067 => x"8d387551",
  1068 => x"abcf2dbd",
  1069 => x"980856a1",
  1070 => x"c7047382",
  1071 => x"d4d52e87",
  1072 => x"38b88051",
  1073 => x"a28904be",
  1074 => x"80527551",
  1075 => x"9cdd2dbd",
  1076 => x"980855bd",
  1077 => x"9808802e",
  1078 => x"83de3888",
  1079 => x"53b7f452",
  1080 => x"bed2519d",
  1081 => x"fd2dbd98",
  1082 => x"088a3881",
  1083 => x"0b80c48c",
  1084 => x"0ca28f04",
  1085 => x"8853b7e8",
  1086 => x"52beb651",
  1087 => x"9dfd2dbd",
  1088 => x"9808802e",
  1089 => x"8a38b894",
  1090 => x"5185fe2d",
  1091 => x"a2eb0480",
  1092 => x"c1fe0b80",
  1093 => x"f52d5473",
  1094 => x"80d52e09",
  1095 => x"810680cb",
  1096 => x"3880c1ff",
  1097 => x"0b80f52d",
  1098 => x"547381aa",
  1099 => x"2e098106",
  1100 => x"ba38800b",
  1101 => x"be800b80",
  1102 => x"f52d5654",
  1103 => x"7481e92e",
  1104 => x"83388154",
  1105 => x"7481eb2e",
  1106 => x"8c388055",
  1107 => x"73752e09",
  1108 => x"810682e4",
  1109 => x"38be8b0b",
  1110 => x"80f52d55",
  1111 => x"748d38be",
  1112 => x"8c0b80f5",
  1113 => x"2d547382",
  1114 => x"2e863880",
  1115 => x"55a5b804",
  1116 => x"be8d0b80",
  1117 => x"f52d7080",
  1118 => x"c4840cff",
  1119 => x"0580c488",
  1120 => x"0cbe8e0b",
  1121 => x"80f52dbe",
  1122 => x"8f0b80f5",
  1123 => x"2d587605",
  1124 => x"77828029",
  1125 => x"057080c4",
  1126 => x"940cbe90",
  1127 => x"0b80f52d",
  1128 => x"7080c4a8",
  1129 => x"0c80c48c",
  1130 => x"08595758",
  1131 => x"76802e81",
  1132 => x"ac388853",
  1133 => x"b7f452be",
  1134 => x"d2519dfd",
  1135 => x"2dbd9808",
  1136 => x"81f63880",
  1137 => x"c4840870",
  1138 => x"842b80c4",
  1139 => x"900c7080",
  1140 => x"c4a40cbe",
  1141 => x"a50b80f5",
  1142 => x"2dbea40b",
  1143 => x"80f52d71",
  1144 => x"82802905",
  1145 => x"bea60b80",
  1146 => x"f52d7084",
  1147 => x"80802912",
  1148 => x"bea70b80",
  1149 => x"f52d7081",
  1150 => x"800a2912",
  1151 => x"7080c4ac",
  1152 => x"0c80c4a8",
  1153 => x"08712980",
  1154 => x"c4940805",
  1155 => x"7080c498",
  1156 => x"0cbead0b",
  1157 => x"80f52dbe",
  1158 => x"ac0b80f5",
  1159 => x"2d718280",
  1160 => x"2905beae",
  1161 => x"0b80f52d",
  1162 => x"70848080",
  1163 => x"2912beaf",
  1164 => x"0b80f52d",
  1165 => x"70982b81",
  1166 => x"f00a0672",
  1167 => x"057080c4",
  1168 => x"9c0cfe11",
  1169 => x"7e297705",
  1170 => x"80c4a00c",
  1171 => x"52595243",
  1172 => x"545e5152",
  1173 => x"59525d57",
  1174 => x"5957a5b1",
  1175 => x"04be920b",
  1176 => x"80f52dbe",
  1177 => x"910b80f5",
  1178 => x"2d718280",
  1179 => x"29057080",
  1180 => x"c4900c70",
  1181 => x"a02983ff",
  1182 => x"0570892a",
  1183 => x"7080c4a4",
  1184 => x"0cbe970b",
  1185 => x"80f52dbe",
  1186 => x"960b80f5",
  1187 => x"2d718280",
  1188 => x"29057080",
  1189 => x"c4ac0c7b",
  1190 => x"71291e70",
  1191 => x"80c4a00c",
  1192 => x"7d80c49c",
  1193 => x"0c730580",
  1194 => x"c4980c55",
  1195 => x"5e515155",
  1196 => x"5580519e",
  1197 => x"bb2d8155",
  1198 => x"74bd980c",
  1199 => x"02a8050d",
  1200 => x"0402ec05",
  1201 => x"0d767087",
  1202 => x"2c7180ff",
  1203 => x"06555654",
  1204 => x"80c48c08",
  1205 => x"8a387388",
  1206 => x"2c7481ff",
  1207 => x"065455be",
  1208 => x"805280c4",
  1209 => x"94081551",
  1210 => x"9cdd2dbd",
  1211 => x"980854bd",
  1212 => x"9808802e",
  1213 => x"b43880c4",
  1214 => x"8c08802e",
  1215 => x"98387284",
  1216 => x"29be8005",
  1217 => x"70085253",
  1218 => x"abcf2dbd",
  1219 => x"9808f00a",
  1220 => x"0653a6a7",
  1221 => x"047210be",
  1222 => x"80057080",
  1223 => x"e02d5253",
  1224 => x"abff2dbd",
  1225 => x"98085372",
  1226 => x"5473bd98",
  1227 => x"0c029405",
  1228 => x"0d0402e0",
  1229 => x"050d7970",
  1230 => x"842c80c4",
  1231 => x"b4080571",
  1232 => x"8f065255",
  1233 => x"53728938",
  1234 => x"be805273",
  1235 => x"519cdd2d",
  1236 => x"72a029be",
  1237 => x"80055480",
  1238 => x"7480f52d",
  1239 => x"56537473",
  1240 => x"2e833881",
  1241 => x"537481e5",
  1242 => x"2e81f138",
  1243 => x"81707406",
  1244 => x"54587280",
  1245 => x"2e81e538",
  1246 => x"8b1480f5",
  1247 => x"2d70832a",
  1248 => x"79065856",
  1249 => x"769938bb",
  1250 => x"dc085372",
  1251 => x"89387280",
  1252 => x"c2800b81",
  1253 => x"b72d76bb",
  1254 => x"dc0c7353",
  1255 => x"a8de0475",
  1256 => x"8f2e0981",
  1257 => x"0681b538",
  1258 => x"749f068d",
  1259 => x"2980c1f3",
  1260 => x"11515381",
  1261 => x"1480f52d",
  1262 => x"73708105",
  1263 => x"5581b72d",
  1264 => x"831480f5",
  1265 => x"2d737081",
  1266 => x"055581b7",
  1267 => x"2d851480",
  1268 => x"f52d7370",
  1269 => x"81055581",
  1270 => x"b72d8714",
  1271 => x"80f52d73",
  1272 => x"70810555",
  1273 => x"81b72d89",
  1274 => x"1480f52d",
  1275 => x"73708105",
  1276 => x"5581b72d",
  1277 => x"8e1480f5",
  1278 => x"2d737081",
  1279 => x"055581b7",
  1280 => x"2d901480",
  1281 => x"f52d7370",
  1282 => x"81055581",
  1283 => x"b72d9214",
  1284 => x"80f52d73",
  1285 => x"70810555",
  1286 => x"81b72d94",
  1287 => x"1480f52d",
  1288 => x"73708105",
  1289 => x"5581b72d",
  1290 => x"961480f5",
  1291 => x"2d737081",
  1292 => x"055581b7",
  1293 => x"2d981480",
  1294 => x"f52d7370",
  1295 => x"81055581",
  1296 => x"b72d9c14",
  1297 => x"80f52d73",
  1298 => x"70810555",
  1299 => x"81b72d9e",
  1300 => x"1480f52d",
  1301 => x"7381b72d",
  1302 => x"77bbdc0c",
  1303 => x"805372bd",
  1304 => x"980c02a0",
  1305 => x"050d0402",
  1306 => x"cc050d7e",
  1307 => x"605e5a80",
  1308 => x"0b80c4b0",
  1309 => x"0880c4b4",
  1310 => x"08595c56",
  1311 => x"805880c4",
  1312 => x"9008782e",
  1313 => x"81b03877",
  1314 => x"8f06a017",
  1315 => x"5754738f",
  1316 => x"38be8052",
  1317 => x"76518117",
  1318 => x"579cdd2d",
  1319 => x"be805680",
  1320 => x"7680f52d",
  1321 => x"56547474",
  1322 => x"2e833881",
  1323 => x"547481e5",
  1324 => x"2e80f738",
  1325 => x"81707506",
  1326 => x"555c7380",
  1327 => x"2e80eb38",
  1328 => x"8b1680f5",
  1329 => x"2d980659",
  1330 => x"7880df38",
  1331 => x"8b537c52",
  1332 => x"75519dfd",
  1333 => x"2dbd9808",
  1334 => x"80d0389c",
  1335 => x"160851ab",
  1336 => x"cf2dbd98",
  1337 => x"08841b0c",
  1338 => x"9a1680e0",
  1339 => x"2d51abff",
  1340 => x"2dbd9808",
  1341 => x"bd980888",
  1342 => x"1c0cbd98",
  1343 => x"08555580",
  1344 => x"c48c0880",
  1345 => x"2e983894",
  1346 => x"1680e02d",
  1347 => x"51abff2d",
  1348 => x"bd980890",
  1349 => x"2b83fff0",
  1350 => x"0a067016",
  1351 => x"51547388",
  1352 => x"1b0c787a",
  1353 => x"0c7b54aa",
  1354 => x"ef048118",
  1355 => x"5880c490",
  1356 => x"087826fe",
  1357 => x"d23880c4",
  1358 => x"8c08802e",
  1359 => x"b0387a51",
  1360 => x"a5c12dbd",
  1361 => x"9808bd98",
  1362 => x"0880ffff",
  1363 => x"fff80655",
  1364 => x"5b7380ff",
  1365 => x"fffff82e",
  1366 => x"9438bd98",
  1367 => x"08fe0580",
  1368 => x"c4840829",
  1369 => x"80c49808",
  1370 => x"0557a8fc",
  1371 => x"04805473",
  1372 => x"bd980c02",
  1373 => x"b4050d04",
  1374 => x"02f4050d",
  1375 => x"74700881",
  1376 => x"05710c70",
  1377 => x"0880c488",
  1378 => x"08065353",
  1379 => x"718e3888",
  1380 => x"130851a5",
  1381 => x"c12dbd98",
  1382 => x"0888140c",
  1383 => x"810bbd98",
  1384 => x"0c028c05",
  1385 => x"0d0402f0",
  1386 => x"050d7588",
  1387 => x"1108fe05",
  1388 => x"80c48408",
  1389 => x"2980c498",
  1390 => x"08117208",
  1391 => x"80c48808",
  1392 => x"06057955",
  1393 => x"5354549c",
  1394 => x"dd2d0290",
  1395 => x"050d0402",
  1396 => x"f4050d74",
  1397 => x"70882a83",
  1398 => x"fe800670",
  1399 => x"72982a07",
  1400 => x"72882b87",
  1401 => x"fc808006",
  1402 => x"73982b81",
  1403 => x"f00a0671",
  1404 => x"730707bd",
  1405 => x"980c5651",
  1406 => x"5351028c",
  1407 => x"050d0402",
  1408 => x"f8050d02",
  1409 => x"8e0580f5",
  1410 => x"2d74882b",
  1411 => x"077083ff",
  1412 => x"ff06bd98",
  1413 => x"0c510288",
  1414 => x"050d0402",
  1415 => x"f4050d74",
  1416 => x"76785354",
  1417 => x"52807125",
  1418 => x"97387270",
  1419 => x"81055480",
  1420 => x"f52d7270",
  1421 => x"81055481",
  1422 => x"b72dff11",
  1423 => x"5170eb38",
  1424 => x"807281b7",
  1425 => x"2d028c05",
  1426 => x"0d0402e8",
  1427 => x"050d7756",
  1428 => x"80705654",
  1429 => x"737624b3",
  1430 => x"3880c490",
  1431 => x"08742eab",
  1432 => x"387351a6",
  1433 => x"b22dbd98",
  1434 => x"08bd9808",
  1435 => x"09810570",
  1436 => x"bd980807",
  1437 => x"9f2a7705",
  1438 => x"81175757",
  1439 => x"53537476",
  1440 => x"24893880",
  1441 => x"c4900874",
  1442 => x"26d73872",
  1443 => x"bd980c02",
  1444 => x"98050d04",
  1445 => x"02f0050d",
  1446 => x"bd940816",
  1447 => x"51acca2d",
  1448 => x"bd980880",
  1449 => x"2e9e388b",
  1450 => x"53bd9808",
  1451 => x"5280c280",
  1452 => x"51ac9b2d",
  1453 => x"80c4bc08",
  1454 => x"5473802e",
  1455 => x"873880c2",
  1456 => x"8051732d",
  1457 => x"0290050d",
  1458 => x"0402dc05",
  1459 => x"0d80705a",
  1460 => x"5574bd94",
  1461 => x"0825b138",
  1462 => x"80c49008",
  1463 => x"752ea938",
  1464 => x"7851a6b2",
  1465 => x"2dbd9808",
  1466 => x"09810570",
  1467 => x"bd980807",
  1468 => x"9f2a7605",
  1469 => x"811b5b56",
  1470 => x"5474bd94",
  1471 => x"08258938",
  1472 => x"80c49008",
  1473 => x"7926d938",
  1474 => x"80557880",
  1475 => x"c4900827",
  1476 => x"81d43878",
  1477 => x"51a6b22d",
  1478 => x"bd980880",
  1479 => x"2e81a838",
  1480 => x"bd98088b",
  1481 => x"0580f52d",
  1482 => x"70842a70",
  1483 => x"81067710",
  1484 => x"78842b80",
  1485 => x"c2800b80",
  1486 => x"f52d5c5c",
  1487 => x"53515556",
  1488 => x"73802e80",
  1489 => x"c9387416",
  1490 => x"822bb08a",
  1491 => x"0bbbe812",
  1492 => x"0c547775",
  1493 => x"311080c4",
  1494 => x"c0115556",
  1495 => x"90747081",
  1496 => x"055681b7",
  1497 => x"2da07481",
  1498 => x"b72d7681",
  1499 => x"ff068116",
  1500 => x"58547380",
  1501 => x"2e8a389c",
  1502 => x"5380c280",
  1503 => x"52af8604",
  1504 => x"8b53bd98",
  1505 => x"085280c4",
  1506 => x"c21651af",
  1507 => x"bf047416",
  1508 => x"822bad94",
  1509 => x"0bbbe812",
  1510 => x"0c547681",
  1511 => x"ff068116",
  1512 => x"58547380",
  1513 => x"2e8a389c",
  1514 => x"5380c280",
  1515 => x"52afb604",
  1516 => x"8b53bd98",
  1517 => x"08527775",
  1518 => x"311080c4",
  1519 => x"c0055176",
  1520 => x"55ac9b2d",
  1521 => x"afdb0474",
  1522 => x"90297531",
  1523 => x"701080c4",
  1524 => x"c0055154",
  1525 => x"bd980874",
  1526 => x"81b72d81",
  1527 => x"1959748b",
  1528 => x"24a338ae",
  1529 => x"8a047490",
  1530 => x"29753170",
  1531 => x"1080c4c0",
  1532 => x"058c7731",
  1533 => x"57515480",
  1534 => x"7481b72d",
  1535 => x"9e14ff16",
  1536 => x"565474f3",
  1537 => x"3802a405",
  1538 => x"0d0402fc",
  1539 => x"050dbd94",
  1540 => x"081351ac",
  1541 => x"ca2dbd98",
  1542 => x"08802e88",
  1543 => x"38bd9808",
  1544 => x"519ebb2d",
  1545 => x"800bbd94",
  1546 => x"0cadc92d",
  1547 => x"8ff22d02",
  1548 => x"84050d04",
  1549 => x"02fc050d",
  1550 => x"725170fd",
  1551 => x"2ead3870",
  1552 => x"fd248a38",
  1553 => x"70fc2e80",
  1554 => x"c438b195",
  1555 => x"0470fe2e",
  1556 => x"b13870ff",
  1557 => x"2e098106",
  1558 => x"bc38bd94",
  1559 => x"08517080",
  1560 => x"2eb338ff",
  1561 => x"11bd940c",
  1562 => x"b19504bd",
  1563 => x"9408f005",
  1564 => x"70bd940c",
  1565 => x"51708025",
  1566 => x"9c38800b",
  1567 => x"bd940cb1",
  1568 => x"9504bd94",
  1569 => x"088105bd",
  1570 => x"940cb195",
  1571 => x"04bd9408",
  1572 => x"9005bd94",
  1573 => x"0cadc92d",
  1574 => x"8ff22d02",
  1575 => x"84050d04",
  1576 => x"02fc050d",
  1577 => x"800bbd94",
  1578 => x"0cadc92d",
  1579 => x"8f892dbd",
  1580 => x"9808bd84",
  1581 => x"0cbbe051",
  1582 => x"918d2d02",
  1583 => x"84050d04",
  1584 => x"7180c4bc",
  1585 => x"0c040000",
  1586 => x"00ffffff",
  1587 => x"ff00ffff",
  1588 => x"ffff00ff",
  1589 => x"ffffff00",
  1590 => x"52657365",
  1591 => x"74000000",
  1592 => x"43617267",
  1593 => x"61722044",
  1594 => x"6973636f",
  1595 => x"2f43696e",
  1596 => x"74612010",
  1597 => x"00000000",
  1598 => x"45786974",
  1599 => x"00000000",
  1600 => x"46444320",
  1601 => x"4f726967",
  1602 => x"696e616c",
  1603 => x"00000000",
  1604 => x"46444320",
  1605 => x"46617374",
  1606 => x"00000000",
  1607 => x"4d756c74",
  1608 => x"69666163",
  1609 => x"65203220",
  1610 => x"456e6162",
  1611 => x"6c656400",
  1612 => x"4d756c74",
  1613 => x"69666163",
  1614 => x"65203220",
  1615 => x"48696464",
  1616 => x"656e0000",
  1617 => x"4d756c74",
  1618 => x"69666163",
  1619 => x"65203220",
  1620 => x"44697361",
  1621 => x"626c6564",
  1622 => x"00000000",
  1623 => x"4d6f7573",
  1624 => x"65204469",
  1625 => x"7361626c",
  1626 => x"65640000",
  1627 => x"4d6f7573",
  1628 => x"6520456e",
  1629 => x"61626c65",
  1630 => x"64000000",
  1631 => x"506c6179",
  1632 => x"63697479",
  1633 => x"20446973",
  1634 => x"61626c65",
  1635 => x"64000000",
  1636 => x"506c6179",
  1637 => x"63697479",
  1638 => x"20456e61",
  1639 => x"626c6564",
  1640 => x"00000000",
  1641 => x"52696768",
  1642 => x"74205368",
  1643 => x"69667420",
  1644 => x"61732042",
  1645 => x"61636b73",
  1646 => x"6c617368",
  1647 => x"00000000",
  1648 => x"52696768",
  1649 => x"74205368",
  1650 => x"69667420",
  1651 => x"61732053",
  1652 => x"68696674",
  1653 => x"00000000",
  1654 => x"536f756e",
  1655 => x"64206f75",
  1656 => x"74707574",
  1657 => x"20537465",
  1658 => x"72656f00",
  1659 => x"536f756e",
  1660 => x"64206f75",
  1661 => x"74707574",
  1662 => x"204d6f6e",
  1663 => x"6f000000",
  1664 => x"54617065",
  1665 => x"20736f75",
  1666 => x"6e642044",
  1667 => x"69736162",
  1668 => x"6c656400",
  1669 => x"54617065",
  1670 => x"20736f75",
  1671 => x"6e642045",
  1672 => x"6e61626c",
  1673 => x"65640000",
  1674 => x"43505520",
  1675 => x"74696d69",
  1676 => x"6e677320",
  1677 => x"4f726967",
  1678 => x"696e616c",
  1679 => x"00000000",
  1680 => x"43505520",
  1681 => x"74696d69",
  1682 => x"6e677320",
  1683 => x"46617374",
  1684 => x"00000000",
  1685 => x"53696e63",
  1686 => x"20736967",
  1687 => x"6e616c73",
  1688 => x"204f7269",
  1689 => x"67696e61",
  1690 => x"6c000000",
  1691 => x"53696e63",
  1692 => x"20736967",
  1693 => x"6e616c73",
  1694 => x"2046696c",
  1695 => x"74657265",
  1696 => x"64000000",
  1697 => x"43525443",
  1698 => x"20547970",
  1699 => x"65203100",
  1700 => x"43525443",
  1701 => x"20547970",
  1702 => x"65203200",
  1703 => x"44697370",
  1704 => x"6c617920",
  1705 => x"436f6c6f",
  1706 => x"72284741",
  1707 => x"29000000",
  1708 => x"44697370",
  1709 => x"6c617920",
  1710 => x"436f6c6f",
  1711 => x"72202841",
  1712 => x"53494329",
  1713 => x"00000000",
  1714 => x"44697370",
  1715 => x"6c617920",
  1716 => x"47726565",
  1717 => x"6e000000",
  1718 => x"44697370",
  1719 => x"6c617920",
  1720 => x"416d6265",
  1721 => x"72000000",
  1722 => x"44697370",
  1723 => x"6c617920",
  1724 => x"4379616e",
  1725 => x"00000000",
  1726 => x"44697370",
  1727 => x"6c617920",
  1728 => x"57686974",
  1729 => x"65000000",
  1730 => x"5363616e",
  1731 => x"6c696e65",
  1732 => x"73204e6f",
  1733 => x"6e650000",
  1734 => x"5363616e",
  1735 => x"6c696e65",
  1736 => x"73204352",
  1737 => x"54203235",
  1738 => x"25000000",
  1739 => x"5363616e",
  1740 => x"6c696e65",
  1741 => x"73204352",
  1742 => x"54203530",
  1743 => x"25000000",
  1744 => x"5363616e",
  1745 => x"6c696e65",
  1746 => x"73204352",
  1747 => x"54203735",
  1748 => x"25000000",
  1749 => x"43617267",
  1750 => x"61204661",
  1751 => x"6c6c6964",
  1752 => x"61000000",
  1753 => x"4f4b0000",
  1754 => x"414d5354",
  1755 => x"52414420",
  1756 => x"44415400",
  1757 => x"16200000",
  1758 => x"14200000",
  1759 => x"15200000",
  1760 => x"53442069",
  1761 => x"6e69742e",
  1762 => x"2e2e0a00",
  1763 => x"53442063",
  1764 => x"61726420",
  1765 => x"72657365",
  1766 => x"74206661",
  1767 => x"696c6564",
  1768 => x"210a0000",
  1769 => x"53444843",
  1770 => x"20657272",
  1771 => x"6f72210a",
  1772 => x"00000000",
  1773 => x"57726974",
  1774 => x"65206661",
  1775 => x"696c6564",
  1776 => x"0a000000",
  1777 => x"52656164",
  1778 => x"20666169",
  1779 => x"6c65640a",
  1780 => x"00000000",
  1781 => x"43617264",
  1782 => x"20696e69",
  1783 => x"74206661",
  1784 => x"696c6564",
  1785 => x"0a000000",
  1786 => x"46415431",
  1787 => x"36202020",
  1788 => x"00000000",
  1789 => x"46415433",
  1790 => x"32202020",
  1791 => x"00000000",
  1792 => x"4e6f2070",
  1793 => x"61727469",
  1794 => x"74696f6e",
  1795 => x"20736967",
  1796 => x"0a000000",
  1797 => x"42616420",
  1798 => x"70617274",
  1799 => x"0a000000",
  1800 => x"4261636b",
  1801 => x"00000000",
  1802 => x"00000002",
  1803 => x"00000002",
  1804 => x"000018d8",
  1805 => x"0000034e",
  1806 => x"00000003",
  1807 => x"00001d58",
  1808 => x"00000004",
  1809 => x"00000003",
  1810 => x"00001d40",
  1811 => x"00000006",
  1812 => x"00000003",
  1813 => x"00001d38",
  1814 => x"00000002",
  1815 => x"00000003",
  1816 => x"00001d30",
  1817 => x"00000002",
  1818 => x"00000003",
  1819 => x"00001d28",
  1820 => x"00000002",
  1821 => x"00000003",
  1822 => x"00001d20",
  1823 => x"00000002",
  1824 => x"00000003",
  1825 => x"00001d18",
  1826 => x"00000002",
  1827 => x"00000003",
  1828 => x"00001d10",
  1829 => x"00000002",
  1830 => x"00000003",
  1831 => x"00001d08",
  1832 => x"00000002",
  1833 => x"00000003",
  1834 => x"00001d00",
  1835 => x"00000002",
  1836 => x"00000003",
  1837 => x"00001cf4",
  1838 => x"00000003",
  1839 => x"00000003",
  1840 => x"00001cec",
  1841 => x"00000002",
  1842 => x"00000002",
  1843 => x"000018e0",
  1844 => x"000018a0",
  1845 => x"00000002",
  1846 => x"000018f8",
  1847 => x"00000790",
  1848 => x"00000000",
  1849 => x"00000000",
  1850 => x"00000000",
  1851 => x"00001900",
  1852 => x"00001910",
  1853 => x"0000191c",
  1854 => x"00001930",
  1855 => x"00001944",
  1856 => x"0000195c",
  1857 => x"0000196c",
  1858 => x"0000197c",
  1859 => x"00001990",
  1860 => x"000019a4",
  1861 => x"000019c0",
  1862 => x"000019d8",
  1863 => x"000019ec",
  1864 => x"00001a00",
  1865 => x"00001a14",
  1866 => x"00001a28",
  1867 => x"00001a40",
  1868 => x"00001a54",
  1869 => x"00001a6c",
  1870 => x"00001a84",
  1871 => x"00001a90",
  1872 => x"00001a9c",
  1873 => x"00001ab0",
  1874 => x"00001ac8",
  1875 => x"00001ad8",
  1876 => x"00001ae8",
  1877 => x"00001af8",
  1878 => x"00001b08",
  1879 => x"00001b18",
  1880 => x"00001b2c",
  1881 => x"00001b40",
  1882 => x"00000004",
  1883 => x"00001b54",
  1884 => x"00001d68",
  1885 => x"00000004",
  1886 => x"00001b64",
  1887 => x"00001c2c",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"00000000",
  1895 => x"00000000",
  1896 => x"00000000",
  1897 => x"00000000",
  1898 => x"00000000",
  1899 => x"00000000",
  1900 => x"00000000",
  1901 => x"00000000",
  1902 => x"00000000",
  1903 => x"00000000",
  1904 => x"00000000",
  1905 => x"00000000",
  1906 => x"00000000",
  1907 => x"00000000",
  1908 => x"00000000",
  1909 => x"00000000",
  1910 => x"00000000",
  1911 => x"00000000",
  1912 => x"00000002",
  1913 => x"00002240",
  1914 => x"00001694",
  1915 => x"00000002",
  1916 => x"0000225e",
  1917 => x"00001694",
  1918 => x"00000002",
  1919 => x"0000227c",
  1920 => x"00001694",
  1921 => x"00000002",
  1922 => x"0000229a",
  1923 => x"00001694",
  1924 => x"00000002",
  1925 => x"000022b8",
  1926 => x"00001694",
  1927 => x"00000002",
  1928 => x"000022d6",
  1929 => x"00001694",
  1930 => x"00000002",
  1931 => x"000022f4",
  1932 => x"00001694",
  1933 => x"00000002",
  1934 => x"00002312",
  1935 => x"00001694",
  1936 => x"00000002",
  1937 => x"00002330",
  1938 => x"00001694",
  1939 => x"00000002",
  1940 => x"0000234e",
  1941 => x"00001694",
  1942 => x"00000002",
  1943 => x"0000236c",
  1944 => x"00001694",
  1945 => x"00000002",
  1946 => x"0000238a",
  1947 => x"00001694",
  1948 => x"00000002",
  1949 => x"000023a8",
  1950 => x"00001694",
  1951 => x"00000004",
  1952 => x"00001c20",
  1953 => x"00000000",
  1954 => x"00000000",
  1955 => x"00000000",
  1956 => x"00001834",
  1957 => x"00000000",
	others => x"00000000"
);

begin

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memAWriteEnable = '1') and (from_zpu.memBWriteEnable = '1') and (from_zpu.memAAddr=from_zpu.memBAddr) and (from_zpu.memAWrite/=from_zpu.memBWrite) then
			report "write collision" severity failure;
		end if;
	
		if (from_zpu.memAWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memAWrite;
			to_zpu.memARead <= from_zpu.memAWrite;
		else
			to_zpu.memARead <= ram(to_integer(unsigned(from_zpu.memAAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;

process (clk)
begin
	if (clk'event and clk = '1') then
		if (from_zpu.memBWriteEnable = '1') then
			ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2)))) := from_zpu.memBWrite;
			to_zpu.memBRead <= from_zpu.memBWrite;
		else
			to_zpu.memBRead <= ram(to_integer(unsigned(from_zpu.memBAddr(maxAddrBitBRAM downto 2))));
		end if;
	end if;
end process;


end arch;

